`timescale 1ns/100ps
module gf128mul(
    input       [6:0] a,
    input       [6:0] b,
    output  reg [6:0] z
);
always @(*)
begin
    case (b)
        7'd1:
            begin
                z[0] = a[0];
                z[1] = a[1];
                z[2] = a[2];
                z[3] = a[3];
                z[4] = a[4];
                z[5] = a[5];
                z[6] = a[6];
            end
        7'd4:
            begin
                z[0] = a[5];
                z[1] = a[6];
                z[2] = a[0];
                z[3] = a[1] ^ a[5];
                z[4] = a[2] ^ a[6];
                z[5] = a[3];
                z[6] = a[4];
            end
        7'd6:
            begin
                z[0] = a[5] ^ a[6];
                z[1] = a[0] ^ a[6];
                z[2] = a[0] ^ a[1];
                z[3] = a[1] ^ a[2] ^ a[5] ^ a[6];
                z[4] = a[2] ^ a[3] ^ a[6];
                z[5] = a[3] ^ a[4];
                z[6] = a[4] ^ a[5];
            end
        7'd8:
            begin
                z[0] = a[4];
                z[1] = a[5];
                z[2] = a[6];
                z[3] = a[0] ^ a[4];
                z[4] = a[1] ^ a[5];
                z[5] = a[2] ^ a[6];
                z[6] = a[3];
            end
        7'd10:
            begin
                z[0] = a[4] ^ a[6];
                z[1] = a[0] ^ a[5];
                z[2] = a[1] ^ a[6];
                z[3] = a[0] ^ a[2] ^ a[4] ^ a[6];
                z[4] = a[1] ^ a[3] ^ a[5];
                z[5] = a[2] ^ a[4] ^ a[6];
                z[6] = a[3] ^ a[5];
            end
        7'd15:
            begin
                z[0] = a[0] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[3] ^ a[4] ^ a[5] ^ a[6];
            end
        7'd20:
            begin
                z[0] = a[3] ^ a[5];
                z[1] = a[4] ^ a[6];
                z[2] = a[0] ^ a[5];
                z[3] = a[1] ^ a[3] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[2] ^ a[4] ^ a[6];
                z[5] = a[1] ^ a[3] ^ a[5];
                z[6] = a[2] ^ a[4] ^ a[6];
            end
        7'd21:
            begin
                z[0] = a[0] ^ a[3] ^ a[5];
                z[1] = a[1] ^ a[4] ^ a[6];
                z[2] = a[0] ^ a[2] ^ a[5];
                z[3] = a[1] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[2] ^ a[6];
                z[5] = a[1] ^ a[3];
                z[6] = a[2] ^ a[4];
            end
        7'd24:
            begin
                z[0] = a[3] ^ a[4];
                z[1] = a[4] ^ a[5];
                z[2] = a[5] ^ a[6];
                z[3] = a[0] ^ a[3] ^ a[4] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[4] ^ a[5];
                z[5] = a[1] ^ a[2] ^ a[5] ^ a[6];
                z[6] = a[2] ^ a[3] ^ a[6];
            end
        7'd26:
            begin
                z[0] = a[3] ^ a[4] ^ a[6];
                z[1] = a[0] ^ a[4] ^ a[5];
                z[2] = a[1] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5];
                z[5] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[2] ^ a[3] ^ a[5] ^ a[6];
            end
        7'd27:
            begin
                z[0] = a[0] ^ a[3] ^ a[4] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[4] ^ a[5];
                z[2] = a[1] ^ a[2] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[2] ^ a[4];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[5];
                z[5] = a[1] ^ a[2] ^ a[4] ^ a[6];
                z[6] = a[2] ^ a[3] ^ a[5];
            end
        7'd30:
            begin
                z[0] = a[3] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[0] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
            end
        7'd32:
            begin
                z[0] = a[2] ^ a[6];
                z[1] = a[3];
                z[2] = a[4];
                z[3] = a[2] ^ a[5] ^ a[6];
                z[4] = a[3] ^ a[6];
                z[5] = a[0] ^ a[4];
                z[6] = a[1] ^ a[5];
            end
        7'd35:
            begin
                z[0] = a[0] ^ a[2];
                z[1] = a[0] ^ a[1] ^ a[3];
                z[2] = a[1] ^ a[2] ^ a[4];
                z[3] = a[3] ^ a[5];
                z[4] = a[4] ^ a[6];
                z[5] = a[0] ^ a[5];
                z[6] = a[1] ^ a[6];
            end
        7'd36:
            begin
                z[0] = a[2] ^ a[5] ^ a[6];
                z[1] = a[3] ^ a[6];
                z[2] = a[0] ^ a[4];
                z[3] = a[1] ^ a[2] ^ a[6];
                z[4] = a[2] ^ a[3];
                z[5] = a[0] ^ a[3] ^ a[4];
                z[6] = a[1] ^ a[4] ^ a[5];
            end
        7'd37:
            begin
                z[0] = a[0] ^ a[2] ^ a[5] ^ a[6];
                z[1] = a[1] ^ a[3] ^ a[6];
                z[2] = a[0] ^ a[2] ^ a[4];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[6];
                z[4] = a[2] ^ a[3] ^ a[4];
                z[5] = a[0] ^ a[3] ^ a[4] ^ a[5];
                z[6] = a[1] ^ a[4] ^ a[5] ^ a[6];
            end
        7'd39:
            begin
                z[0] = a[0] ^ a[2] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[4];
                z[3] = a[1] ^ a[3];
                z[4] = a[2] ^ a[4];
                z[5] = a[0] ^ a[3] ^ a[5];
                z[6] = a[1] ^ a[4] ^ a[6];
            end
        7'd49:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[6];
                z[1] = a[1] ^ a[3] ^ a[4];
                z[2] = a[2] ^ a[4] ^ a[5];
                z[3] = a[2] ^ a[5];
                z[4] = a[0] ^ a[3] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[4];
                z[6] = a[1] ^ a[2] ^ a[5];
            end
        7'd50:
            begin
                z[0] = a[2] ^ a[3];
                z[1] = a[0] ^ a[3] ^ a[4];
                z[2] = a[1] ^ a[4] ^ a[5];
                z[3] = a[3] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[4] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[5];
                z[6] = a[1] ^ a[2] ^ a[6];
            end
        7'd52:
            begin
                z[0] = a[2] ^ a[3] ^ a[5] ^ a[6];
                z[1] = a[3] ^ a[4] ^ a[6];
                z[2] = a[0] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[2] ^ a[3];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5];
                z[6] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
            end
        7'd55:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[6];
                z[4] = a[0] ^ a[2];
                z[5] = a[0] ^ a[1] ^ a[3];
                z[6] = a[1] ^ a[2] ^ a[4];
            end
        7'd58:
            begin
                z[0] = a[2] ^ a[3] ^ a[4];
                z[1] = a[0] ^ a[3] ^ a[4] ^ a[5];
                z[2] = a[1] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[6];
            end
        7'd60:
            begin
                z[0] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[3] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
            end
        7'd62:
            begin
                z[0] = a[2] ^ a[3] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
            end
        7'd63:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[4] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[5];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[4];
            end
        7'd64:
            begin
                z[0] = a[1] ^ a[5];
                z[1] = a[2] ^ a[6];
                z[2] = a[3];
                z[3] = a[1] ^ a[4] ^ a[5];
                z[4] = a[2] ^ a[5] ^ a[6];
                z[5] = a[3] ^ a[6];
                z[6] = a[0] ^ a[4];
            end
        7'd65:
            begin
                z[0] = a[0] ^ a[1] ^ a[5];
                z[1] = a[1] ^ a[2] ^ a[6];
                z[2] = a[2] ^ a[3];
                z[3] = a[1] ^ a[3] ^ a[4] ^ a[5];
                z[4] = a[2] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[3] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[4] ^ a[6];
            end
        7'd70:
            begin
                z[0] = a[1] ^ a[6];
                z[1] = a[0] ^ a[2];
                z[2] = a[0] ^ a[1] ^ a[3];
                z[3] = a[2] ^ a[4] ^ a[6];
                z[4] = a[3] ^ a[5];
                z[5] = a[4] ^ a[6];
                z[6] = a[0] ^ a[5];
            end
        7'd72:
            begin
                z[0] = a[1] ^ a[4] ^ a[5];
                z[1] = a[2] ^ a[5] ^ a[6];
                z[2] = a[3] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[5];
                z[4] = a[1] ^ a[2] ^ a[6];
                z[5] = a[2] ^ a[3];
                z[6] = a[0] ^ a[3] ^ a[4];
            end
        7'd76:
            begin
                z[0] = a[1] ^ a[4];
                z[1] = a[2] ^ a[5];
                z[2] = a[0] ^ a[3] ^ a[6];
                z[3] = a[0];
                z[4] = a[1];
                z[5] = a[2];
                z[6] = a[0] ^ a[3];
            end
        7'd77:
            begin
                z[0] = a[0] ^ a[1] ^ a[4];
                z[1] = a[1] ^ a[2] ^ a[5];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[6];
                z[3] = a[0] ^ a[3];
                z[4] = a[1] ^ a[4];
                z[5] = a[2] ^ a[5];
                z[6] = a[0] ^ a[3] ^ a[6];
            end
        7'd79:
            begin
                z[0] = a[0] ^ a[1] ^ a[4] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[5];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[6];
                z[4] = a[1] ^ a[3] ^ a[4];
                z[5] = a[2] ^ a[4] ^ a[5];
                z[6] = a[0] ^ a[3] ^ a[5] ^ a[6];
            end
        7'd80:
            begin
                z[0] = a[1] ^ a[3] ^ a[5];
                z[1] = a[2] ^ a[4] ^ a[6];
                z[2] = a[3] ^ a[5];
                z[3] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[1] ^ a[3] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[2] ^ a[4] ^ a[6];
            end
        7'd81:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[5];
                z[1] = a[1] ^ a[2] ^ a[4] ^ a[6];
                z[2] = a[2] ^ a[3] ^ a[5];
                z[3] = a[1] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[2] ^ a[5] ^ a[6];
                z[5] = a[1] ^ a[3] ^ a[6];
                z[6] = a[0] ^ a[2] ^ a[4];
            end
        7'd87:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[4];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5];
                z[3] = a[2] ^ a[4];
                z[4] = a[0] ^ a[3] ^ a[5];
                z[5] = a[1] ^ a[4] ^ a[6];
                z[6] = a[0] ^ a[2] ^ a[5];
            end
        7'd89:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5];
                z[1] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[2] ^ a[3] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[6];
                z[5] = a[1] ^ a[2] ^ a[3];
                z[6] = a[0] ^ a[2] ^ a[3] ^ a[4];
            end
        7'd92:
            begin
                z[0] = a[1] ^ a[3] ^ a[4];
                z[1] = a[2] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[3] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[3] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[4];
                z[5] = a[1] ^ a[2] ^ a[5];
                z[6] = a[0] ^ a[2] ^ a[3] ^ a[6];
            end
        7'd96:
            begin
                z[0] = a[1] ^ a[2] ^ a[5] ^ a[6];
                z[1] = a[2] ^ a[3] ^ a[6];
                z[2] = a[3] ^ a[4];
                z[3] = a[1] ^ a[2] ^ a[4] ^ a[6];
                z[4] = a[2] ^ a[3] ^ a[5];
                z[5] = a[0] ^ a[3] ^ a[4] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[4] ^ a[5];
            end
        7'd97:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[6];
                z[2] = a[2] ^ a[3] ^ a[4];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[4] = a[2] ^ a[3] ^ a[4] ^ a[5];
                z[5] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6];
            end
        7'd101:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[6];
                z[1] = a[1] ^ a[2] ^ a[3];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[3] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[3] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[5] ^ a[6];
            end
        7'd103:
            begin
                z[0] = a[0] ^ a[1] ^ a[2];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
                z[3] = a[3] ^ a[4] ^ a[5];
                z[4] = a[4] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[6];
            end
        7'd104:
            begin
                z[0] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[2] ^ a[3] ^ a[5] ^ a[6];
                z[2] = a[3] ^ a[4] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[6];
                z[4] = a[1] ^ a[2] ^ a[3];
                z[5] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[6] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5];
            end
        7'd108:
            begin
                z[0] = a[1] ^ a[2] ^ a[4] ^ a[6];
                z[1] = a[2] ^ a[3] ^ a[5];
                z[2] = a[0] ^ a[3] ^ a[4] ^ a[6];
                z[3] = a[0] ^ a[2] ^ a[5] ^ a[6];
                z[4] = a[1] ^ a[3] ^ a[6];
                z[5] = a[0] ^ a[2] ^ a[4];
                z[6] = a[0] ^ a[1] ^ a[3] ^ a[5];
            end
        7'd114:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[5];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[2] = a[1] ^ a[3] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[3] ^ a[4] ^ a[6];
                z[4] = a[0] ^ a[2] ^ a[4] ^ a[5];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[6];
            end
        7'd116:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[6];
                z[1] = a[2] ^ a[3] ^ a[4];
                z[2] = a[0] ^ a[3] ^ a[4] ^ a[5];
                z[3] = a[2] ^ a[3] ^ a[4] ^ a[5];
                z[4] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6];
            end
        7'd118:
            begin
                z[0] = a[1] ^ a[2] ^ a[3];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5];
                z[3] = a[3] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[6];
            end
        7'd120:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[3] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
            end
        7'd122:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[4];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
            end
        7'd124:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[1] = a[2] ^ a[3] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[5];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
            end
        7'd125:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[2] ^ a[5];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[4];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5];
            end
        7'd126:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[4];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[3] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[4] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[5];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6];
            end
        7'd127:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[2];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3];
            end
        default:
            begin
                z[0] = 0; 
                z[1] = 0; 
                z[2] = 0; 
                z[3] = 0; 
                z[4] = 0; 
                z[5] = 0; 
                z[6] = 0; 
            end
    endcase
end
endmodule
