`timescale 1ns/100ps
module gf64mul(
    input       [5:0] a,
    input       [5:0] b,
    output  reg [5:0] z
);
always @(*)
begin
    case (b)
        6'd1:
            begin
                z[0] = a[0];
                z[1] = a[1];
                z[2] = a[2];
                z[3] = a[3];
                z[4] = a[4];
                z[5] = a[5];
            end
        6'd2:
            begin
                z[0] = a[5];
                z[1] = a[0] ^ a[5];
                z[2] = a[1];
                z[3] = a[2];
                z[4] = a[3];
                z[5] = a[4];
            end
        6'd4:
            begin
                z[0] = a[4];
                z[1] = a[4] ^ a[5];
                z[2] = a[0] ^ a[5];
                z[3] = a[1];
                z[4] = a[2];
                z[5] = a[3];
            end
        6'd5:
            begin
                z[0] = a[0] ^ a[4];
                z[1] = a[1] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[2] ^ a[5];
                z[3] = a[1] ^ a[3];
                z[4] = a[2] ^ a[4];
                z[5] = a[3] ^ a[5];
            end
        6'd6:
            begin
                z[0] = a[4] ^ a[5];
                z[1] = a[0] ^ a[4];
                z[2] = a[0] ^ a[1] ^ a[5];
                z[3] = a[1] ^ a[2];
                z[4] = a[2] ^ a[3];
                z[5] = a[3] ^ a[4];
            end
        6'd8:
            begin
                z[0] = a[3];
                z[1] = a[3] ^ a[4];
                z[2] = a[4] ^ a[5];
                z[3] = a[0] ^ a[5];
                z[4] = a[1];
                z[5] = a[2];
            end
        6'd10:
            begin
                z[0] = a[3] ^ a[5];
                z[1] = a[0] ^ a[3] ^ a[4] ^ a[5];
                z[2] = a[1] ^ a[4] ^ a[5];
                z[3] = a[0] ^ a[2] ^ a[5];
                z[4] = a[1] ^ a[3];
                z[5] = a[2] ^ a[4];
            end
        6'd12:
            begin
                z[0] = a[3] ^ a[4];
                z[1] = a[3] ^ a[5];
                z[2] = a[0] ^ a[4];
                z[3] = a[0] ^ a[1] ^ a[5];
                z[4] = a[1] ^ a[2];
                z[5] = a[2] ^ a[3];
            end
        6'd13:
            begin
                z[0] = a[0] ^ a[3] ^ a[4];
                z[1] = a[1] ^ a[3] ^ a[5];
                z[2] = a[0] ^ a[2] ^ a[4];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[5];
                z[4] = a[1] ^ a[2] ^ a[4];
                z[5] = a[2] ^ a[3] ^ a[5];
            end
        6'd14:
            begin
                z[0] = a[3] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[3];
                z[2] = a[0] ^ a[1] ^ a[4];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[5];
                z[4] = a[1] ^ a[2] ^ a[3];
                z[5] = a[2] ^ a[3] ^ a[4];
            end
        6'd17:
            begin
                z[0] = a[0] ^ a[2];
                z[1] = a[1] ^ a[2] ^ a[3];
                z[2] = a[2] ^ a[3] ^ a[4];
                z[3] = a[3] ^ a[4] ^ a[5];
                z[4] = a[0] ^ a[4] ^ a[5];
                z[5] = a[1] ^ a[5];
            end
        6'd18:
            begin
                z[0] = a[2] ^ a[5];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[5];
                z[2] = a[1] ^ a[3] ^ a[4];
                z[3] = a[2] ^ a[4] ^ a[5];
                z[4] = a[0] ^ a[3] ^ a[5];
                z[5] = a[1] ^ a[4];
            end
        6'd19:
            begin
                z[0] = a[0] ^ a[2] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5];
                z[2] = a[1] ^ a[2] ^ a[3] ^ a[4];
                z[3] = a[2] ^ a[3] ^ a[4] ^ a[5];
                z[4] = a[0] ^ a[3] ^ a[4] ^ a[5];
                z[5] = a[1] ^ a[4] ^ a[5];
            end
        6'd20:
            begin
                z[0] = a[2] ^ a[4];
                z[1] = a[2] ^ a[3] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[3] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[4] ^ a[5];
                z[4] = a[0] ^ a[2] ^ a[5];
                z[5] = a[1] ^ a[3];
            end
        6'd21:
            begin
                z[0] = a[0] ^ a[2] ^ a[4];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[3] ^ a[4] ^ a[5];
                z[4] = a[0] ^ a[2] ^ a[4] ^ a[5];
                z[5] = a[1] ^ a[3] ^ a[5];
            end
        6'd22:
            begin
                z[0] = a[2] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[2] ^ a[4] ^ a[5];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[5];
                z[5] = a[1] ^ a[3] ^ a[4];
            end
        6'd23:
            begin
                z[0] = a[0] ^ a[2] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[5] = a[1] ^ a[3] ^ a[4] ^ a[5];
            end
        6'd25:
            begin
                z[0] = a[0] ^ a[2] ^ a[3];
                z[1] = a[1] ^ a[2] ^ a[4];
                z[2] = a[2] ^ a[3] ^ a[5];
                z[3] = a[0] ^ a[3] ^ a[4];
                z[4] = a[0] ^ a[1] ^ a[4] ^ a[5];
                z[5] = a[1] ^ a[2] ^ a[5];
            end
        6'd26:
            begin
                z[0] = a[2] ^ a[3] ^ a[5];
                z[1] = a[0] ^ a[2] ^ a[4] ^ a[5];
                z[2] = a[1] ^ a[3] ^ a[5];
                z[3] = a[0] ^ a[2] ^ a[4];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[5];
                z[5] = a[1] ^ a[2] ^ a[4];
            end
        6'd27:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5];
                z[2] = a[1] ^ a[2] ^ a[3] ^ a[5];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5];
                z[5] = a[1] ^ a[2] ^ a[4] ^ a[5];
            end
        6'd28:
            begin
                z[0] = a[2] ^ a[3] ^ a[4];
                z[1] = a[2] ^ a[5];
                z[2] = a[0] ^ a[3];
                z[3] = a[0] ^ a[1] ^ a[4];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[5];
                z[5] = a[1] ^ a[2] ^ a[3];
            end
        6'd29:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[1] = a[1] ^ a[2] ^ a[5];
                z[2] = a[0] ^ a[2] ^ a[3];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[4];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[5];
            end
        6'd30:
            begin
                z[0] = a[2] ^ a[3] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[2];
                z[2] = a[0] ^ a[1] ^ a[3];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[4];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[4];
            end
        6'd31:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[2];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
            end
        6'd34:
            begin
                z[0] = a[1] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[5];
                z[2] = a[1] ^ a[2] ^ a[3];
                z[3] = a[2] ^ a[3] ^ a[4];
                z[4] = a[3] ^ a[4] ^ a[5];
                z[5] = a[0] ^ a[4] ^ a[5];
            end
        6'd35:
            begin
                z[0] = a[0] ^ a[1] ^ a[5];
                z[1] = a[0] ^ a[2] ^ a[5];
                z[2] = a[1] ^ a[3];
                z[3] = a[2] ^ a[4];
                z[4] = a[3] ^ a[5];
                z[5] = a[0] ^ a[4];
            end
        6'd36:
            begin
                z[0] = a[1] ^ a[4];
                z[1] = a[1] ^ a[2] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[5];
                z[3] = a[1] ^ a[3] ^ a[4];
                z[4] = a[2] ^ a[4] ^ a[5];
                z[5] = a[0] ^ a[3] ^ a[5];
            end
        6'd37:
            begin
                z[0] = a[0] ^ a[1] ^ a[4];
                z[1] = a[2] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[3] ^ a[5];
                z[3] = a[1] ^ a[4];
                z[4] = a[2] ^ a[5];
                z[5] = a[0] ^ a[3];
            end
        6'd38:
            begin
                z[0] = a[1] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[4];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[4];
                z[4] = a[2] ^ a[3] ^ a[4] ^ a[5];
                z[5] = a[0] ^ a[3] ^ a[4] ^ a[5];
            end
        6'd41:
            begin
                z[0] = a[0] ^ a[1] ^ a[3];
                z[1] = a[2] ^ a[3] ^ a[4];
                z[2] = a[3] ^ a[4] ^ a[5];
                z[3] = a[0] ^ a[4] ^ a[5];
                z[4] = a[1] ^ a[5];
                z[5] = a[0] ^ a[2];
            end
        6'd46:
            begin
                z[0] = a[1] ^ a[3] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[5] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
            end
        6'd47:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[2] ^ a[3];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[4];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[5];
                z[5] = a[0] ^ a[2] ^ a[3] ^ a[4];
            end
        6'd48:
            begin
                z[0] = a[1] ^ a[2];
                z[1] = a[1] ^ a[3];
                z[2] = a[2] ^ a[4];
                z[3] = a[3] ^ a[5];
                z[4] = a[0] ^ a[4];
                z[5] = a[0] ^ a[1] ^ a[5];
            end
        6'd49:
            begin
                z[0] = a[0] ^ a[1] ^ a[2];
                z[1] = a[3];
                z[2] = a[4];
                z[3] = a[5];
                z[4] = a[0];
                z[5] = a[0] ^ a[1];
            end
        6'd50:
            begin
                z[0] = a[1] ^ a[2] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[5];
                z[2] = a[1] ^ a[2] ^ a[4];
                z[3] = a[2] ^ a[3] ^ a[5];
                z[4] = a[0] ^ a[3] ^ a[4];
                z[5] = a[0] ^ a[1] ^ a[4] ^ a[5];
            end
        6'd52:
            begin
                z[0] = a[1] ^ a[2] ^ a[4];
                z[1] = a[1] ^ a[3] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[2] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[3] ^ a[5];
                z[4] = a[0] ^ a[2] ^ a[4];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[5];
            end
        6'd53:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[4];
                z[1] = a[3] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[5];
                z[4] = a[0] ^ a[2];
                z[5] = a[0] ^ a[1] ^ a[3];
            end
        6'd54:
            begin
                z[0] = a[1] ^ a[2] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[4];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[5];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5];
            end
        6'd55:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[3] ^ a[4];
                z[2] = a[0] ^ a[1] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[2] ^ a[5];
                z[4] = a[0] ^ a[2] ^ a[3];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[4];
            end
        6'd57:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3];
                z[1] = a[4];
                z[2] = a[5];
                z[3] = a[0];
                z[4] = a[0] ^ a[1];
                z[5] = a[0] ^ a[1] ^ a[2];
            end
        6'd59:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5];
                z[1] = a[0] ^ a[4] ^ a[5];
                z[2] = a[1] ^ a[5];
                z[3] = a[0] ^ a[2];
                z[4] = a[0] ^ a[1] ^ a[3];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[4];
            end
        6'd61:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
                z[1] = a[5];
                z[2] = a[0];
                z[3] = a[0] ^ a[1];
                z[4] = a[0] ^ a[1] ^ a[2];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3];
            end
        6'd62:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[1];
                z[2] = a[0] ^ a[1] ^ a[2];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
            end
        default:
            begin
                z[0] = 0; 
                z[1] = 0; 
                z[2] = 0; 
                z[3] = 0; 
                z[4] = 0; 
                z[5] = 0; 
            end
    endcase
end
endmodule
