`define BLK_NUM    2
`define SYM_BW    4
`define N_NUM    15
`define R_NUM    4
