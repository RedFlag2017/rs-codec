`timescale 1ns/100ps
module gf256mul_dec(
    input       [7:0] a,
    input       [7:0] b,
    output  reg [7:0] z
);
always @(*)
begin
    case (b)
        8'd1:
            begin
                z[0] = a[0];
                z[1] = a[1];
                z[2] = a[2];
                z[3] = a[3];
                z[4] = a[4];
                z[5] = a[5];
                z[6] = a[6];
                z[7] = a[7];
            end
        8'd2:
            begin
                z[0] = a[7];
                z[1] = a[0];
                z[2] = a[1] ^ a[7];
                z[3] = a[2] ^ a[7];
                z[4] = a[3] ^ a[7];
                z[5] = a[4];
                z[6] = a[5];
                z[7] = a[6];
            end
        8'd3:
            begin
                z[0] = a[0] ^ a[7];
                z[1] = a[0] ^ a[1];
                z[2] = a[1] ^ a[2] ^ a[7];
                z[3] = a[2] ^ a[3] ^ a[7];
                z[4] = a[3] ^ a[4] ^ a[7];
                z[5] = a[4] ^ a[5];
                z[6] = a[5] ^ a[6];
                z[7] = a[6] ^ a[7];
            end
        8'd4:
            begin
                z[0] = a[6];
                z[1] = a[7];
                z[2] = a[0] ^ a[6];
                z[3] = a[1] ^ a[6] ^ a[7];
                z[4] = a[2] ^ a[6] ^ a[7];
                z[5] = a[3] ^ a[7];
                z[6] = a[4];
                z[7] = a[5];
            end
        8'd5:
            begin
                z[0] = a[0] ^ a[6];
                z[1] = a[1] ^ a[7];
                z[2] = a[0] ^ a[2] ^ a[6];
                z[3] = a[1] ^ a[3] ^ a[6] ^ a[7];
                z[4] = a[2] ^ a[4] ^ a[6] ^ a[7];
                z[5] = a[3] ^ a[5] ^ a[7];
                z[6] = a[4] ^ a[6];
                z[7] = a[5] ^ a[7];
            end
        8'd6:
            begin
                z[0] = a[6] ^ a[7];
                z[1] = a[0] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[6] ^ a[7];
                z[3] = a[1] ^ a[2] ^ a[6];
                z[4] = a[2] ^ a[3] ^ a[6];
                z[5] = a[3] ^ a[4] ^ a[7];
                z[6] = a[4] ^ a[5];
                z[7] = a[5] ^ a[6];
            end
        8'd7:
            begin
                z[0] = a[0] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[6] ^ a[7];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[6];
                z[4] = a[2] ^ a[3] ^ a[4] ^ a[6];
                z[5] = a[3] ^ a[4] ^ a[5] ^ a[7];
                z[6] = a[4] ^ a[5] ^ a[6];
                z[7] = a[5] ^ a[6] ^ a[7];
            end
        8'd8:
            begin
                z[0] = a[5];
                z[1] = a[6];
                z[2] = a[5] ^ a[7];
                z[3] = a[0] ^ a[5] ^ a[6];
                z[4] = a[1] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[2] ^ a[6] ^ a[7];
                z[6] = a[3] ^ a[7];
                z[7] = a[4];
            end
        8'd9:
            begin
                z[0] = a[0] ^ a[5];
                z[1] = a[1] ^ a[6];
                z[2] = a[2] ^ a[5] ^ a[7];
                z[3] = a[0] ^ a[3] ^ a[5] ^ a[6];
                z[4] = a[1] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[2] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[3] ^ a[6] ^ a[7];
                z[7] = a[4] ^ a[7];
            end
        8'd10:
            begin
                z[0] = a[5] ^ a[7];
                z[1] = a[0] ^ a[6];
                z[2] = a[1] ^ a[5];
                z[3] = a[0] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[1] ^ a[3] ^ a[5] ^ a[6];
                z[5] = a[2] ^ a[4] ^ a[6] ^ a[7];
                z[6] = a[3] ^ a[5] ^ a[7];
                z[7] = a[4] ^ a[6];
            end
        8'd11:
            begin
                z[0] = a[0] ^ a[5] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[6];
                z[2] = a[1] ^ a[2] ^ a[5];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[3] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[4] ^ a[6] ^ a[7];
            end
        8'd12:
            begin
                z[0] = a[5] ^ a[6];
                z[1] = a[6] ^ a[7];
                z[2] = a[0] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[5] ^ a[7];
                z[4] = a[1] ^ a[2] ^ a[5];
                z[5] = a[2] ^ a[3] ^ a[6];
                z[6] = a[3] ^ a[4] ^ a[7];
                z[7] = a[4] ^ a[5];
            end
        8'd13:
            begin
                z[0] = a[0] ^ a[5] ^ a[6];
                z[1] = a[1] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[7];
                z[4] = a[1] ^ a[2] ^ a[4] ^ a[5];
                z[5] = a[2] ^ a[3] ^ a[5] ^ a[6];
                z[6] = a[3] ^ a[4] ^ a[6] ^ a[7];
                z[7] = a[4] ^ a[5] ^ a[7];
            end
        8'd14:
            begin
                z[0] = a[5] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[5];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[5] = a[2] ^ a[3] ^ a[4] ^ a[6];
                z[6] = a[3] ^ a[4] ^ a[5] ^ a[7];
                z[7] = a[4] ^ a[5] ^ a[6];
            end
        8'd15:
            begin
                z[0] = a[0] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[5] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[4] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd16:
            begin
                z[0] = a[4];
                z[1] = a[5];
                z[2] = a[4] ^ a[6];
                z[3] = a[4] ^ a[5] ^ a[7];
                z[4] = a[0] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[1] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[2] ^ a[6] ^ a[7];
                z[7] = a[3] ^ a[7];
            end
        8'd17:
            begin
                z[0] = a[0] ^ a[4];
                z[1] = a[1] ^ a[5];
                z[2] = a[2] ^ a[4] ^ a[6];
                z[3] = a[3] ^ a[4] ^ a[5] ^ a[7];
                z[4] = a[0] ^ a[5] ^ a[6];
                z[5] = a[1] ^ a[6] ^ a[7];
                z[6] = a[2] ^ a[7];
                z[7] = a[3];
            end
        8'd18:
            begin
                z[0] = a[4] ^ a[7];
                z[1] = a[0] ^ a[5];
                z[2] = a[1] ^ a[4] ^ a[6] ^ a[7];
                z[3] = a[2] ^ a[4] ^ a[5];
                z[4] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[1] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[2] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[3] ^ a[6] ^ a[7];
            end
        8'd19:
            begin
                z[0] = a[0] ^ a[4] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[5];
                z[2] = a[1] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[3] = a[2] ^ a[3] ^ a[4] ^ a[5];
                z[4] = a[0] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[1] ^ a[4] ^ a[6] ^ a[7];
                z[6] = a[2] ^ a[5] ^ a[7];
                z[7] = a[3] ^ a[6];
            end
        8'd20:
            begin
                z[0] = a[4] ^ a[6];
                z[1] = a[5] ^ a[7];
                z[2] = a[0] ^ a[4];
                z[3] = a[1] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[5] = a[1] ^ a[3] ^ a[5] ^ a[6];
                z[6] = a[2] ^ a[4] ^ a[6] ^ a[7];
                z[7] = a[3] ^ a[5] ^ a[7];
            end
        8'd21:
            begin
                z[0] = a[0] ^ a[4] ^ a[6];
                z[1] = a[1] ^ a[5] ^ a[7];
                z[2] = a[0] ^ a[2] ^ a[4];
                z[3] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[2] ^ a[5] ^ a[7];
                z[5] = a[1] ^ a[3] ^ a[6];
                z[6] = a[2] ^ a[4] ^ a[7];
                z[7] = a[3] ^ a[5];
            end
        8'd22:
            begin
                z[0] = a[4] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[5] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[4] ^ a[7];
                z[3] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[5] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[3] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd23:
            begin
                z[0] = a[0] ^ a[4] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[5] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[7];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[5];
                z[5] = a[1] ^ a[3] ^ a[4] ^ a[6];
                z[6] = a[2] ^ a[4] ^ a[5] ^ a[7];
                z[7] = a[3] ^ a[5] ^ a[6];
            end
        8'd24:
            begin
                z[0] = a[4] ^ a[5];
                z[1] = a[5] ^ a[6];
                z[2] = a[4] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[4] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[4] ^ a[7];
                z[5] = a[1] ^ a[2] ^ a[5];
                z[6] = a[2] ^ a[3] ^ a[6];
                z[7] = a[3] ^ a[4] ^ a[7];
            end
        8'd25:
            begin
                z[0] = a[0] ^ a[4] ^ a[5];
                z[1] = a[1] ^ a[5] ^ a[6];
                z[2] = a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[7];
                z[5] = a[1] ^ a[2];
                z[6] = a[2] ^ a[3];
                z[7] = a[3] ^ a[4];
            end
        8'd26:
            begin
                z[0] = a[4] ^ a[5] ^ a[7];
                z[1] = a[0] ^ a[5] ^ a[6];
                z[2] = a[1] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[2] ^ a[4] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[4];
                z[5] = a[1] ^ a[2] ^ a[4] ^ a[5];
                z[6] = a[2] ^ a[3] ^ a[5] ^ a[6];
                z[7] = a[3] ^ a[4] ^ a[6] ^ a[7];
            end
        8'd27:
            begin
                z[0] = a[0] ^ a[4] ^ a[5] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[5] ^ a[6];
                z[2] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[3];
                z[5] = a[1] ^ a[2] ^ a[4];
                z[6] = a[2] ^ a[3] ^ a[5];
                z[7] = a[3] ^ a[4] ^ a[6];
            end
        8'd28:
            begin
                z[0] = a[4] ^ a[5] ^ a[6];
                z[1] = a[5] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[4] ^ a[5] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[4];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[6];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[6] = a[2] ^ a[3] ^ a[4] ^ a[6];
                z[7] = a[3] ^ a[4] ^ a[5] ^ a[7];
            end
        8'd29:
            begin
                z[0] = a[0] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[1] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[4];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[6];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[7];
                z[6] = a[2] ^ a[3] ^ a[4];
                z[7] = a[3] ^ a[4] ^ a[5];
            end
        8'd30:
            begin
                z[0] = a[4] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[4] ^ a[5];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[6] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[7] = a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd31:
            begin
                z[0] = a[0] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[6] = a[2] ^ a[3] ^ a[4] ^ a[5];
                z[7] = a[3] ^ a[4] ^ a[5] ^ a[6];
            end
        8'd32:
            begin
                z[0] = a[3] ^ a[7];
                z[1] = a[4];
                z[2] = a[3] ^ a[5] ^ a[7];
                z[3] = a[3] ^ a[4] ^ a[6] ^ a[7];
                z[4] = a[3] ^ a[4] ^ a[5];
                z[5] = a[0] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[1] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[2] ^ a[6] ^ a[7];
            end
        8'd33:
            begin
                z[0] = a[0] ^ a[3] ^ a[7];
                z[1] = a[1] ^ a[4];
                z[2] = a[2] ^ a[3] ^ a[5] ^ a[7];
                z[3] = a[4] ^ a[6] ^ a[7];
                z[4] = a[3] ^ a[5];
                z[5] = a[0] ^ a[4] ^ a[6];
                z[6] = a[1] ^ a[5] ^ a[7];
                z[7] = a[2] ^ a[6];
            end
        8'd34:
            begin
                z[0] = a[3];
                z[1] = a[0] ^ a[4];
                z[2] = a[1] ^ a[3] ^ a[5];
                z[3] = a[2] ^ a[3] ^ a[4] ^ a[6];
                z[4] = a[4] ^ a[5] ^ a[7];
                z[5] = a[0] ^ a[5] ^ a[6];
                z[6] = a[1] ^ a[6] ^ a[7];
                z[7] = a[2] ^ a[7];
            end
        8'd35:
            begin
                z[0] = a[0] ^ a[3];
                z[1] = a[0] ^ a[1] ^ a[4];
                z[2] = a[1] ^ a[2] ^ a[3] ^ a[5];
                z[3] = a[2] ^ a[4] ^ a[6];
                z[4] = a[5] ^ a[7];
                z[5] = a[0] ^ a[6];
                z[6] = a[1] ^ a[7];
                z[7] = a[2];
            end
        8'd36:
            begin
                z[0] = a[3] ^ a[6] ^ a[7];
                z[1] = a[4] ^ a[7];
                z[2] = a[0] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[1] ^ a[3] ^ a[4];
                z[4] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[1] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[2] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd37:
            begin
                z[0] = a[0] ^ a[3] ^ a[6] ^ a[7];
                z[1] = a[1] ^ a[4] ^ a[7];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[1] ^ a[4];
                z[4] = a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[6] = a[1] ^ a[4] ^ a[5] ^ a[7];
                z[7] = a[2] ^ a[5] ^ a[6];
            end
        8'd38:
            begin
                z[0] = a[3] ^ a[6];
                z[1] = a[0] ^ a[4] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[6];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[4] = a[2] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[1] ^ a[4] ^ a[6] ^ a[7];
                z[7] = a[2] ^ a[5] ^ a[7];
            end
        8'd39:
            begin
                z[0] = a[0] ^ a[3] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[4] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[3] = a[1] ^ a[2] ^ a[4] ^ a[7];
                z[4] = a[2] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[3] ^ a[6] ^ a[7];
                z[6] = a[1] ^ a[4] ^ a[7];
                z[7] = a[2] ^ a[5];
            end
        8'd40:
            begin
                z[0] = a[3] ^ a[5] ^ a[7];
                z[1] = a[4] ^ a[6];
                z[2] = a[3];
                z[3] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[4] = a[1] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[6] = a[1] ^ a[3] ^ a[5] ^ a[6];
                z[7] = a[2] ^ a[4] ^ a[6] ^ a[7];
            end
        8'd41:
            begin
                z[0] = a[0] ^ a[3] ^ a[5] ^ a[7];
                z[1] = a[1] ^ a[4] ^ a[6];
                z[2] = a[2] ^ a[3];
                z[3] = a[0] ^ a[4] ^ a[5] ^ a[7];
                z[4] = a[1] ^ a[3] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[2] ^ a[4] ^ a[7];
                z[6] = a[1] ^ a[3] ^ a[5];
                z[7] = a[2] ^ a[4] ^ a[6];
            end
        8'd42:
            begin
                z[0] = a[3] ^ a[5];
                z[1] = a[0] ^ a[4] ^ a[6];
                z[2] = a[1] ^ a[3] ^ a[7];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[4] = a[1] ^ a[4] ^ a[6];
                z[5] = a[0] ^ a[2] ^ a[5] ^ a[7];
                z[6] = a[1] ^ a[3] ^ a[6];
                z[7] = a[2] ^ a[4] ^ a[7];
            end
        8'd43:
            begin
                z[0] = a[0] ^ a[3] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[4] ^ a[6];
                z[2] = a[1] ^ a[2] ^ a[3] ^ a[7];
                z[3] = a[0] ^ a[2] ^ a[4] ^ a[5];
                z[4] = a[1] ^ a[6];
                z[5] = a[0] ^ a[2] ^ a[7];
                z[6] = a[1] ^ a[3];
                z[7] = a[2] ^ a[4];
            end
        8'd44:
            begin
                z[0] = a[3] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[4] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[3] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[4];
                z[5] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[6] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[7] = a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd45:
            begin
                z[0] = a[0] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[1] ^ a[4] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[1] ^ a[2] ^ a[3];
                z[5] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[6] = a[1] ^ a[3] ^ a[4] ^ a[5];
                z[7] = a[2] ^ a[4] ^ a[5] ^ a[6];
            end
        8'd46:
            begin
                z[0] = a[3] ^ a[5] ^ a[6];
                z[1] = a[0] ^ a[4] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[1] ^ a[2] ^ a[4] ^ a[7];
                z[5] = a[0] ^ a[2] ^ a[3] ^ a[5];
                z[6] = a[1] ^ a[3] ^ a[4] ^ a[6];
                z[7] = a[2] ^ a[4] ^ a[5] ^ a[7];
            end
        8'd47:
            begin
                z[0] = a[0] ^ a[3] ^ a[5] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[4] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[1] ^ a[2] ^ a[7];
                z[5] = a[0] ^ a[2] ^ a[3];
                z[6] = a[1] ^ a[3] ^ a[4];
                z[7] = a[2] ^ a[4] ^ a[5];
            end
        8'd48:
            begin
                z[0] = a[3] ^ a[4] ^ a[7];
                z[1] = a[4] ^ a[5];
                z[2] = a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[3] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[3] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[4] ^ a[7];
                z[6] = a[1] ^ a[2] ^ a[5];
                z[7] = a[2] ^ a[3] ^ a[6];
            end
        8'd49:
            begin
                z[0] = a[0] ^ a[3] ^ a[4] ^ a[7];
                z[1] = a[1] ^ a[4] ^ a[5];
                z[2] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[5] ^ a[6];
                z[4] = a[0] ^ a[3] ^ a[4] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[7];
                z[6] = a[1] ^ a[2] ^ a[5] ^ a[6];
                z[7] = a[2] ^ a[3] ^ a[6] ^ a[7];
            end
        8'd50:
            begin
                z[0] = a[3] ^ a[4];
                z[1] = a[0] ^ a[4] ^ a[5];
                z[2] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[7];
                z[6] = a[1] ^ a[2];
                z[7] = a[2] ^ a[3];
            end
        8'd51:
            begin
                z[0] = a[0] ^ a[3] ^ a[4];
                z[1] = a[0] ^ a[1] ^ a[4] ^ a[5];
                z[2] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[2] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[4] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[5] ^ a[7];
                z[6] = a[1] ^ a[2] ^ a[6];
                z[7] = a[2] ^ a[3] ^ a[7];
            end
        8'd52:
            begin
                z[0] = a[3] ^ a[4] ^ a[6] ^ a[7];
                z[1] = a[4] ^ a[5] ^ a[7];
                z[2] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[3] = a[1] ^ a[3] ^ a[5] ^ a[7];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[4];
                z[6] = a[1] ^ a[2] ^ a[4] ^ a[5];
                z[7] = a[2] ^ a[3] ^ a[5] ^ a[6];
            end
        8'd53:
            begin
                z[0] = a[0] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[1] = a[1] ^ a[4] ^ a[5] ^ a[7];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[3] = a[1] ^ a[5] ^ a[7];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5];
                z[6] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[7] = a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd54:
            begin
                z[0] = a[3] ^ a[4] ^ a[6];
                z[1] = a[0] ^ a[4] ^ a[5] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[5];
                z[4] = a[0] ^ a[2];
                z[5] = a[0] ^ a[1] ^ a[3];
                z[6] = a[1] ^ a[2] ^ a[4];
                z[7] = a[2] ^ a[3] ^ a[5];
            end
        8'd55:
            begin
                z[0] = a[0] ^ a[3] ^ a[4] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[2] ^ a[5];
                z[4] = a[0] ^ a[2] ^ a[4];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[5];
                z[6] = a[1] ^ a[2] ^ a[4] ^ a[6];
                z[7] = a[2] ^ a[3] ^ a[5] ^ a[7];
            end
        8'd56:
            begin
                z[0] = a[3] ^ a[4] ^ a[5] ^ a[7];
                z[1] = a[4] ^ a[5] ^ a[6];
                z[2] = a[3] ^ a[4] ^ a[6];
                z[3] = a[0] ^ a[3];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[6];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[7] = a[2] ^ a[3] ^ a[4] ^ a[6];
            end
        8'd57:
            begin
                z[0] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[1] = a[1] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[2] ^ a[3] ^ a[4] ^ a[6];
                z[3] = a[0];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
            end
        8'd58:
            begin
                z[0] = a[3] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[1] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[5];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[6];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[7];
                z[7] = a[2] ^ a[3] ^ a[4];
            end
        8'd59:
            begin
                z[0] = a[0] ^ a[3] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[2] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[4] ^ a[5];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[7] = a[2] ^ a[3] ^ a[4] ^ a[7];
            end
        8'd60:
            begin
                z[0] = a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[4] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[3] ^ a[4];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[7] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
            end
        8'd61:
            begin
                z[0] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[1] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[3] = a[0] ^ a[1] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd62:
            begin
                z[0] = a[3] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[0] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[7] = a[2] ^ a[3] ^ a[4] ^ a[5];
            end
        8'd63:
            begin
                z[0] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[7] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
            end
        8'd64:
            begin
                z[0] = a[2] ^ a[6] ^ a[7];
                z[1] = a[3] ^ a[7];
                z[2] = a[2] ^ a[4] ^ a[6] ^ a[7];
                z[3] = a[2] ^ a[3] ^ a[5] ^ a[6];
                z[4] = a[2] ^ a[3] ^ a[4];
                z[5] = a[3] ^ a[4] ^ a[5];
                z[6] = a[0] ^ a[4] ^ a[5] ^ a[6];
                z[7] = a[1] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd65:
            begin
                z[0] = a[0] ^ a[2] ^ a[6] ^ a[7];
                z[1] = a[1] ^ a[3] ^ a[7];
                z[2] = a[4] ^ a[6] ^ a[7];
                z[3] = a[2] ^ a[5] ^ a[6];
                z[4] = a[2] ^ a[3];
                z[5] = a[3] ^ a[4];
                z[6] = a[0] ^ a[4] ^ a[5];
                z[7] = a[1] ^ a[5] ^ a[6];
            end
        8'd66:
            begin
                z[0] = a[2] ^ a[6];
                z[1] = a[0] ^ a[3] ^ a[7];
                z[2] = a[1] ^ a[2] ^ a[4] ^ a[6];
                z[3] = a[3] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[2] ^ a[4] ^ a[7];
                z[5] = a[3] ^ a[5];
                z[6] = a[0] ^ a[4] ^ a[6];
                z[7] = a[1] ^ a[5] ^ a[7];
            end
        8'd67:
            begin
                z[0] = a[0] ^ a[2] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[7];
                z[2] = a[1] ^ a[4] ^ a[6];
                z[3] = a[5] ^ a[6] ^ a[7];
                z[4] = a[2] ^ a[7];
                z[5] = a[3];
                z[6] = a[0] ^ a[4];
                z[7] = a[1] ^ a[5];
            end
        8'd68:
            begin
                z[0] = a[2] ^ a[7];
                z[1] = a[3];
                z[2] = a[0] ^ a[2] ^ a[4] ^ a[7];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[4] = a[3] ^ a[4] ^ a[6] ^ a[7];
                z[5] = a[4] ^ a[5] ^ a[7];
                z[6] = a[0] ^ a[5] ^ a[6];
                z[7] = a[1] ^ a[6] ^ a[7];
            end
        8'd69:
            begin
                z[0] = a[0] ^ a[2] ^ a[7];
                z[1] = a[1] ^ a[3];
                z[2] = a[0] ^ a[4] ^ a[7];
                z[3] = a[1] ^ a[2] ^ a[5] ^ a[7];
                z[4] = a[3] ^ a[6] ^ a[7];
                z[5] = a[4] ^ a[7];
                z[6] = a[0] ^ a[5];
                z[7] = a[1] ^ a[6];
            end
        8'd70:
            begin
                z[0] = a[2];
                z[1] = a[0] ^ a[3];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[4];
                z[3] = a[1] ^ a[3] ^ a[5];
                z[4] = a[4] ^ a[6];
                z[5] = a[5] ^ a[7];
                z[6] = a[0] ^ a[6];
                z[7] = a[1] ^ a[7];
            end
        8'd71:
            begin
                z[0] = a[0] ^ a[2];
                z[1] = a[0] ^ a[1] ^ a[3];
                z[2] = a[0] ^ a[1] ^ a[4];
                z[3] = a[1] ^ a[5];
                z[4] = a[6];
                z[5] = a[7];
                z[6] = a[0];
                z[7] = a[1];
            end
        8'd72:
            begin
                z[0] = a[2] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[3] ^ a[6] ^ a[7];
                z[2] = a[2] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[2] ^ a[3];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[1] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd73:
            begin
                z[0] = a[0] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[1] ^ a[3] ^ a[6] ^ a[7];
                z[2] = a[4] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[2];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[7] = a[1] ^ a[4] ^ a[5] ^ a[6];
            end
        8'd74:
            begin
                z[0] = a[2] ^ a[5] ^ a[6];
                z[1] = a[0] ^ a[3] ^ a[6] ^ a[7];
                z[2] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[3] ^ a[7];
                z[4] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[7] = a[1] ^ a[4] ^ a[5] ^ a[7];
            end
        8'd75:
            begin
                z[0] = a[0] ^ a[2] ^ a[5] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[6] ^ a[7];
                z[2] = a[1] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[7];
                z[4] = a[1] ^ a[2] ^ a[5] ^ a[6];
                z[5] = a[2] ^ a[3] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[3] ^ a[4] ^ a[7];
                z[7] = a[1] ^ a[4] ^ a[5];
            end
        8'd76:
            begin
                z[0] = a[2] ^ a[5] ^ a[7];
                z[1] = a[3] ^ a[6];
                z[2] = a[0] ^ a[2] ^ a[4] ^ a[5];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[4] = a[1] ^ a[3] ^ a[4] ^ a[5];
                z[5] = a[2] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[1] ^ a[4] ^ a[6] ^ a[7];
            end
        8'd77:
            begin
                z[0] = a[0] ^ a[2] ^ a[5] ^ a[7];
                z[1] = a[1] ^ a[3] ^ a[6];
                z[2] = a[0] ^ a[4] ^ a[5];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[6] ^ a[7];
                z[4] = a[1] ^ a[3] ^ a[5];
                z[5] = a[2] ^ a[4] ^ a[6];
                z[6] = a[0] ^ a[3] ^ a[5] ^ a[7];
                z[7] = a[1] ^ a[4] ^ a[6];
            end
        8'd78:
            begin
                z[0] = a[2] ^ a[5];
                z[1] = a[0] ^ a[3] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[6];
                z[4] = a[1] ^ a[4] ^ a[5] ^ a[7];
                z[5] = a[2] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[3] ^ a[6] ^ a[7];
                z[7] = a[1] ^ a[4] ^ a[7];
            end
        8'd79:
            begin
                z[0] = a[0] ^ a[2] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[6];
                z[4] = a[1] ^ a[5] ^ a[7];
                z[5] = a[2] ^ a[6];
                z[6] = a[0] ^ a[3] ^ a[7];
                z[7] = a[1] ^ a[4];
            end
        8'd80:
            begin
                z[0] = a[2] ^ a[4] ^ a[6] ^ a[7];
                z[1] = a[3] ^ a[5] ^ a[7];
                z[2] = a[2] ^ a[7];
                z[3] = a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[5] = a[1] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[7] = a[1] ^ a[3] ^ a[5] ^ a[6];
            end
        8'd81:
            begin
                z[0] = a[0] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[1] = a[1] ^ a[3] ^ a[5] ^ a[7];
                z[2] = a[7];
                z[3] = a[2] ^ a[4] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[1] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd82:
            begin
                z[0] = a[2] ^ a[4] ^ a[6];
                z[1] = a[0] ^ a[3] ^ a[5] ^ a[7];
                z[2] = a[1] ^ a[2];
                z[3] = a[3] ^ a[4] ^ a[6];
                z[4] = a[0] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[1] ^ a[3] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[2] ^ a[4] ^ a[7];
                z[7] = a[1] ^ a[3] ^ a[5];
            end
        8'd83:
            begin
                z[0] = a[0] ^ a[2] ^ a[4] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[7];
                z[2] = a[1];
                z[3] = a[4] ^ a[6];
                z[4] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[1] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[7] = a[1] ^ a[3] ^ a[5] ^ a[7];
            end
        8'd84:
            begin
                z[0] = a[2] ^ a[4] ^ a[7];
                z[1] = a[3] ^ a[5];
                z[2] = a[0] ^ a[2] ^ a[6] ^ a[7];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[4];
                z[4] = a[0] ^ a[3] ^ a[5] ^ a[7];
                z[5] = a[1] ^ a[4] ^ a[6];
                z[6] = a[0] ^ a[2] ^ a[5] ^ a[7];
                z[7] = a[1] ^ a[3] ^ a[6];
            end
        8'd85:
            begin
                z[0] = a[0] ^ a[2] ^ a[4] ^ a[7];
                z[1] = a[1] ^ a[3] ^ a[5];
                z[2] = a[0] ^ a[6] ^ a[7];
                z[3] = a[1] ^ a[2] ^ a[4];
                z[4] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[5] = a[1] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[1] ^ a[3] ^ a[6] ^ a[7];
            end
        8'd86:
            begin
                z[0] = a[2] ^ a[4];
                z[1] = a[0] ^ a[3] ^ a[5];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[6];
                z[3] = a[1] ^ a[3] ^ a[4] ^ a[7];
                z[4] = a[0] ^ a[5];
                z[5] = a[1] ^ a[6];
                z[6] = a[0] ^ a[2] ^ a[7];
                z[7] = a[1] ^ a[3];
            end
        8'd87:
            begin
                z[0] = a[0] ^ a[2] ^ a[4];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[5];
                z[2] = a[0] ^ a[1] ^ a[6];
                z[3] = a[1] ^ a[4] ^ a[7];
                z[4] = a[0] ^ a[4] ^ a[5];
                z[5] = a[1] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[2] ^ a[6] ^ a[7];
                z[7] = a[1] ^ a[3] ^ a[7];
            end
        8'd88:
            begin
                z[0] = a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[3] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[2] ^ a[5];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[7];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[4];
                z[6] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[7] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
            end
        8'd89:
            begin
                z[0] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[1] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[5];
                z[3] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[6] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[7] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd90:
            begin
                z[0] = a[2] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[0] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[1] ^ a[2] ^ a[5] ^ a[7];
                z[3] = a[0] ^ a[3] ^ a[4] ^ a[5];
                z[4] = a[0] ^ a[1] ^ a[2];
                z[5] = a[1] ^ a[2] ^ a[3];
                z[6] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[7] = a[1] ^ a[3] ^ a[4] ^ a[5];
            end
        8'd91:
            begin
                z[0] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[1] ^ a[5] ^ a[7];
                z[3] = a[0] ^ a[4] ^ a[5];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[4];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[5];
                z[6] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[7] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
            end
        8'd92:
            begin
                z[0] = a[2] ^ a[4] ^ a[5] ^ a[7];
                z[1] = a[3] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[2] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[6];
                z[5] = a[1] ^ a[2] ^ a[4] ^ a[7];
                z[6] = a[0] ^ a[2] ^ a[3] ^ a[5];
                z[7] = a[1] ^ a[3] ^ a[4] ^ a[6];
            end
        8'd93:
            begin
                z[0] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[1] = a[1] ^ a[3] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6];
                z[5] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[6] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[7] = a[1] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
            end
        8'd94:
            begin
                z[0] = a[2] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[3] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[6] ^ a[7];
                z[5] = a[1] ^ a[2] ^ a[7];
                z[6] = a[0] ^ a[2] ^ a[3];
                z[7] = a[1] ^ a[3] ^ a[4];
            end
        8'd95:
            begin
                z[0] = a[0] ^ a[2] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[4] ^ a[6] ^ a[7];
                z[5] = a[1] ^ a[2] ^ a[5] ^ a[7];
                z[6] = a[0] ^ a[2] ^ a[3] ^ a[6];
                z[7] = a[1] ^ a[3] ^ a[4] ^ a[7];
            end
        8'd96:
            begin
                z[0] = a[2] ^ a[3] ^ a[6];
                z[1] = a[3] ^ a[4] ^ a[7];
                z[2] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[2] ^ a[4] ^ a[5] ^ a[7];
                z[4] = a[2] ^ a[5];
                z[5] = a[0] ^ a[3] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[4] ^ a[7];
                z[7] = a[1] ^ a[2] ^ a[5];
            end
        8'd97:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[6];
                z[1] = a[1] ^ a[3] ^ a[4] ^ a[7];
                z[2] = a[3] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[4] = a[2] ^ a[4] ^ a[5];
                z[5] = a[0] ^ a[3] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[4] ^ a[6] ^ a[7];
                z[7] = a[1] ^ a[2] ^ a[5] ^ a[7];
            end
        8'd98:
            begin
                z[0] = a[2] ^ a[3] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[3] ^ a[4] ^ a[7];
                z[2] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[4] ^ a[5];
                z[4] = a[2] ^ a[3] ^ a[5] ^ a[7];
                z[5] = a[0] ^ a[3] ^ a[4] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[7];
                z[7] = a[1] ^ a[2] ^ a[5] ^ a[6];
            end
        8'd99:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[7];
                z[2] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[3] ^ a[4] ^ a[5];
                z[4] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[5] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[1] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd100:
            begin
                z[0] = a[2] ^ a[3];
                z[1] = a[3] ^ a[4];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[5] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[7];
                z[7] = a[1] ^ a[2];
            end
        8'd101:
            begin
                z[0] = a[0] ^ a[2] ^ a[3];
                z[1] = a[1] ^ a[3] ^ a[4];
                z[2] = a[0] ^ a[3] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[4] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[6] ^ a[7];
                z[7] = a[1] ^ a[2] ^ a[7];
            end
        8'd102:
            begin
                z[0] = a[2] ^ a[3] ^ a[7];
                z[1] = a[0] ^ a[3] ^ a[4];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[3] = a[1] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[3] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[4] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[5] ^ a[7];
                z[7] = a[1] ^ a[2] ^ a[6];
            end
        8'd103:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[4];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[3] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[3] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[1] ^ a[2] ^ a[6] ^ a[7];
            end
        8'd104:
            begin
                z[0] = a[2] ^ a[3] ^ a[5] ^ a[6];
                z[1] = a[3] ^ a[4] ^ a[6] ^ a[7];
                z[2] = a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[4] = a[1] ^ a[2] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[2] ^ a[3] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[3] ^ a[4];
                z[7] = a[1] ^ a[2] ^ a[4] ^ a[5];
            end
        8'd105:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[1] = a[1] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[2] = a[3] ^ a[4] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[4] = a[1] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6];
                z[7] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
            end
        8'd106:
            begin
                z[0] = a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[2] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[3] = a[0] ^ a[4] ^ a[6];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[6];
                z[5] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5];
                z[7] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
            end
        8'd107:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[2] = a[1] ^ a[3] ^ a[4] ^ a[6];
                z[3] = a[0] ^ a[3] ^ a[4] ^ a[6];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[5] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[7] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd108:
            begin
                z[0] = a[2] ^ a[3] ^ a[5];
                z[1] = a[3] ^ a[4] ^ a[6];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[4];
                z[4] = a[1];
                z[5] = a[0] ^ a[2];
                z[6] = a[0] ^ a[1] ^ a[3];
                z[7] = a[1] ^ a[2] ^ a[4];
            end
        8'd109:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[5];
                z[1] = a[1] ^ a[3] ^ a[4] ^ a[6];
                z[2] = a[0] ^ a[3] ^ a[4] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
                z[4] = a[1] ^ a[4];
                z[5] = a[0] ^ a[2] ^ a[5];
                z[6] = a[0] ^ a[1] ^ a[3] ^ a[6];
                z[7] = a[1] ^ a[2] ^ a[4] ^ a[7];
            end
        8'd110:
            begin
                z[0] = a[2] ^ a[3] ^ a[5] ^ a[7];
                z[1] = a[0] ^ a[3] ^ a[4] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
                z[3] = a[0] ^ a[1] ^ a[4] ^ a[7];
                z[4] = a[1] ^ a[3] ^ a[7];
                z[5] = a[0] ^ a[2] ^ a[4];
                z[6] = a[0] ^ a[1] ^ a[3] ^ a[5];
                z[7] = a[1] ^ a[2] ^ a[4] ^ a[6];
            end
        8'd111:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[4];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[7];
                z[4] = a[1] ^ a[3] ^ a[4] ^ a[7];
                z[5] = a[0] ^ a[2] ^ a[4] ^ a[5];
                z[6] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[6];
                z[7] = a[1] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
            end
        8'd112:
            begin
                z[0] = a[2] ^ a[3] ^ a[4] ^ a[6];
                z[1] = a[3] ^ a[4] ^ a[5] ^ a[7];
                z[2] = a[2] ^ a[3] ^ a[5];
                z[3] = a[2];
                z[4] = a[0] ^ a[2] ^ a[4] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[6];
                z[7] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
            end
        8'd113:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[1] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[2] = a[3] ^ a[5];
                z[3] = a[2] ^ a[3];
                z[4] = a[0] ^ a[2] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[4];
                z[7] = a[1] ^ a[2] ^ a[3] ^ a[5];
            end
        8'd114:
            begin
                z[0] = a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[2] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[3] = a[7];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[7] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd115:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[2] = a[1] ^ a[3] ^ a[5] ^ a[7];
                z[3] = a[3] ^ a[7];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5];
                z[7] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
            end
        8'd116:
            begin
                z[0] = a[2] ^ a[3] ^ a[4];
                z[1] = a[3] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[3] = a[1] ^ a[2] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[4] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[5];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[6];
                z[7] = a[1] ^ a[2] ^ a[3] ^ a[7];
            end
        8'd117:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[1] = a[1] ^ a[3] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[3] ^ a[5] ^ a[6];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[7];
                z[5] = a[0] ^ a[1];
                z[6] = a[0] ^ a[1] ^ a[2];
                z[7] = a[1] ^ a[2] ^ a[3];
            end
        8'd118:
            begin
                z[0] = a[2] ^ a[3] ^ a[4] ^ a[7];
                z[1] = a[0] ^ a[3] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[1] ^ a[6];
                z[4] = a[0] ^ a[3] ^ a[4];
                z[5] = a[0] ^ a[1] ^ a[4] ^ a[5];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6];
                z[7] = a[1] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
            end
        8'd119:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[1] ^ a[3] ^ a[6];
                z[4] = a[0] ^ a[3];
                z[5] = a[0] ^ a[1] ^ a[4];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[5];
                z[7] = a[1] ^ a[2] ^ a[3] ^ a[6];
            end
        8'd120:
            begin
                z[0] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[2] ^ a[3] ^ a[7];
                z[3] = a[0] ^ a[2] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[7] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
            end
        8'd121:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[3] ^ a[7];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[7] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
            end
        8'd122:
            begin
                z[0] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[1] ^ a[2] ^ a[3];
                z[3] = a[0] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd123:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[1] ^ a[3];
                z[3] = a[0] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[7] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
            end
        8'd124:
            begin
                z[0] = a[2] ^ a[3] ^ a[4] ^ a[5];
                z[1] = a[3] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[7] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
            end
        8'd125:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[1] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[3] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[7];
                z[7] = a[1] ^ a[2] ^ a[3] ^ a[4];
            end
        8'd126:
            begin
                z[0] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[1] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[5];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
            end
        8'd127:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[5];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[7] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
            end
        8'd128:
            begin
                z[0] = a[1] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[2] ^ a[6] ^ a[7];
                z[2] = a[1] ^ a[3] ^ a[5] ^ a[6];
                z[3] = a[1] ^ a[2] ^ a[4] ^ a[5];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[7];
                z[5] = a[2] ^ a[3] ^ a[4];
                z[6] = a[3] ^ a[4] ^ a[5];
                z[7] = a[0] ^ a[4] ^ a[5] ^ a[6];
            end
        8'd129:
            begin
                z[0] = a[0] ^ a[1] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[1] ^ a[2] ^ a[6] ^ a[7];
                z[2] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[5] = a[2] ^ a[3] ^ a[4] ^ a[5];
                z[6] = a[3] ^ a[4] ^ a[5] ^ a[6];
                z[7] = a[0] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd130:
            begin
                z[0] = a[1] ^ a[5] ^ a[6];
                z[1] = a[0] ^ a[2] ^ a[6] ^ a[7];
                z[2] = a[3] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[1] ^ a[4] ^ a[5] ^ a[7];
                z[4] = a[1] ^ a[2];
                z[5] = a[2] ^ a[3];
                z[6] = a[3] ^ a[4];
                z[7] = a[0] ^ a[4] ^ a[5];
            end
        8'd131:
            begin
                z[0] = a[0] ^ a[1] ^ a[5] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[6] ^ a[7];
                z[2] = a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[4] = a[1] ^ a[2] ^ a[4];
                z[5] = a[2] ^ a[3] ^ a[5];
                z[6] = a[3] ^ a[4] ^ a[6];
                z[7] = a[0] ^ a[4] ^ a[5] ^ a[7];
            end
        8'd132:
            begin
                z[0] = a[1] ^ a[5] ^ a[7];
                z[1] = a[2] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[5];
                z[3] = a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[1] ^ a[3] ^ a[6];
                z[5] = a[2] ^ a[4] ^ a[7];
                z[6] = a[3] ^ a[5];
                z[7] = a[0] ^ a[4] ^ a[6];
            end
        8'd133:
            begin
                z[0] = a[0] ^ a[1] ^ a[5] ^ a[7];
                z[1] = a[1] ^ a[2] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5];
                z[3] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[1] ^ a[3] ^ a[4] ^ a[6];
                z[5] = a[2] ^ a[4] ^ a[5] ^ a[7];
                z[6] = a[3] ^ a[5] ^ a[6];
                z[7] = a[0] ^ a[4] ^ a[6] ^ a[7];
            end
        8'd134:
            begin
                z[0] = a[1] ^ a[5];
                z[1] = a[0] ^ a[2] ^ a[6];
                z[2] = a[0] ^ a[3] ^ a[5] ^ a[7];
                z[3] = a[4] ^ a[5] ^ a[6];
                z[4] = a[1] ^ a[6] ^ a[7];
                z[5] = a[2] ^ a[7];
                z[6] = a[3];
                z[7] = a[0] ^ a[4];
            end
        8'd135:
            begin
                z[0] = a[0] ^ a[1] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[6];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[3] = a[3] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[1] ^ a[4] ^ a[6] ^ a[7];
                z[5] = a[2] ^ a[5] ^ a[7];
                z[6] = a[3] ^ a[6];
                z[7] = a[0] ^ a[4] ^ a[7];
            end
        8'd136:
            begin
                z[0] = a[1] ^ a[6] ^ a[7];
                z[1] = a[2] ^ a[7];
                z[2] = a[1] ^ a[3] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[6];
                z[4] = a[2] ^ a[3] ^ a[5] ^ a[6];
                z[5] = a[3] ^ a[4] ^ a[6] ^ a[7];
                z[6] = a[4] ^ a[5] ^ a[7];
                z[7] = a[0] ^ a[5] ^ a[6];
            end
        8'd137:
            begin
                z[0] = a[0] ^ a[1] ^ a[6] ^ a[7];
                z[1] = a[1] ^ a[2] ^ a[7];
                z[2] = a[1] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[4] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[4] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd138:
            begin
                z[0] = a[1] ^ a[6];
                z[1] = a[0] ^ a[2] ^ a[7];
                z[2] = a[3] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[4] ^ a[6] ^ a[7];
                z[4] = a[2] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[3] ^ a[6] ^ a[7];
                z[6] = a[4] ^ a[7];
                z[7] = a[0] ^ a[5];
            end
        8'd139:
            begin
                z[0] = a[0] ^ a[1] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[7];
                z[2] = a[2] ^ a[3] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[4] = a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[3] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[4] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[5] ^ a[7];
            end
        8'd140:
            begin
                z[0] = a[1] ^ a[7];
                z[1] = a[2];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[7];
                z[3] = a[0] ^ a[2] ^ a[4] ^ a[7];
                z[4] = a[3] ^ a[5] ^ a[7];
                z[5] = a[4] ^ a[6];
                z[6] = a[5] ^ a[7];
                z[7] = a[0] ^ a[6];
            end
        8'd141:
            begin
                z[0] = a[0] ^ a[1] ^ a[7];
                z[1] = a[1] ^ a[2];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[7];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[4] = a[3] ^ a[4] ^ a[5] ^ a[7];
                z[5] = a[4] ^ a[5] ^ a[6];
                z[6] = a[5] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[6] ^ a[7];
            end
        8'd142:
            begin
                z[0] = a[1];
                z[1] = a[0] ^ a[2];
                z[2] = a[0] ^ a[3];
                z[3] = a[0] ^ a[4];
                z[4] = a[5];
                z[5] = a[6];
                z[6] = a[7];
                z[7] = a[0];
            end
        8'd143:
            begin
                z[0] = a[0] ^ a[1];
                z[1] = a[0] ^ a[1] ^ a[2];
                z[2] = a[0] ^ a[2] ^ a[3];
                z[3] = a[0] ^ a[3] ^ a[4];
                z[4] = a[4] ^ a[5];
                z[5] = a[5] ^ a[6];
                z[6] = a[6] ^ a[7];
                z[7] = a[0] ^ a[7];
            end
        8'd144:
            begin
                z[0] = a[1] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[2] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[1] ^ a[3] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[2] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd145:
            begin
                z[0] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[1] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[6] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[7] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
            end
        8'd146:
            begin
                z[0] = a[1] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[0] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[3] ^ a[4] ^ a[5] ^ a[7];
                z[3] = a[1];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
            end
        8'd147:
            begin
                z[0] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[3] = a[1] ^ a[3];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[6] = a[2] ^ a[3] ^ a[4] ^ a[7];
                z[7] = a[0] ^ a[3] ^ a[4] ^ a[5];
            end
        8'd148:
            begin
                z[0] = a[1] ^ a[4] ^ a[5] ^ a[7];
                z[1] = a[2] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[2] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5];
                z[5] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
            end
        8'd149:
            begin
                z[0] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[7];
                z[1] = a[1] ^ a[2] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[2] ^ a[3] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[5];
                z[5] = a[1] ^ a[2] ^ a[4] ^ a[6];
                z[6] = a[2] ^ a[3] ^ a[5] ^ a[7];
                z[7] = a[0] ^ a[3] ^ a[4] ^ a[6];
            end
        8'd150:
            begin
                z[0] = a[1] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[2] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[6] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[7];
                z[5] = a[1] ^ a[2] ^ a[5] ^ a[6];
                z[6] = a[2] ^ a[3] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[3] ^ a[4] ^ a[7];
            end
        8'd151:
            begin
                z[0] = a[0] ^ a[1] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[3] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[5] ^ a[7];
                z[5] = a[1] ^ a[2] ^ a[6];
                z[6] = a[2] ^ a[3] ^ a[7];
                z[7] = a[0] ^ a[3] ^ a[4];
            end
        8'd152:
            begin
                z[0] = a[1] ^ a[4] ^ a[6] ^ a[7];
                z[1] = a[2] ^ a[5] ^ a[7];
                z[2] = a[1] ^ a[3] ^ a[4] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[5] = a[1] ^ a[3] ^ a[4] ^ a[5];
                z[6] = a[2] ^ a[4] ^ a[5] ^ a[6];
                z[7] = a[0] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd153:
            begin
                z[0] = a[0] ^ a[1] ^ a[4] ^ a[6] ^ a[7];
                z[1] = a[1] ^ a[2] ^ a[5] ^ a[7];
                z[2] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[2] ^ a[3];
                z[5] = a[1] ^ a[3] ^ a[4];
                z[6] = a[2] ^ a[4] ^ a[5];
                z[7] = a[0] ^ a[3] ^ a[5] ^ a[6];
            end
        8'd154:
            begin
                z[0] = a[1] ^ a[4] ^ a[6];
                z[1] = a[0] ^ a[2] ^ a[5] ^ a[7];
                z[2] = a[3] ^ a[4];
                z[3] = a[0] ^ a[1] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[2] ^ a[4] ^ a[7];
                z[5] = a[1] ^ a[3] ^ a[5];
                z[6] = a[2] ^ a[4] ^ a[6];
                z[7] = a[0] ^ a[3] ^ a[5] ^ a[7];
            end
        8'd155:
            begin
                z[0] = a[0] ^ a[1] ^ a[4] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[7];
                z[2] = a[2] ^ a[3] ^ a[4];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[2] ^ a[7];
                z[5] = a[1] ^ a[3];
                z[6] = a[2] ^ a[4];
                z[7] = a[0] ^ a[3] ^ a[5];
            end
        8'd156:
            begin
                z[0] = a[1] ^ a[4] ^ a[7];
                z[1] = a[2] ^ a[5];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[2] ^ a[5];
                z[4] = a[0] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[5] = a[1] ^ a[4] ^ a[5] ^ a[7];
                z[6] = a[2] ^ a[5] ^ a[6];
                z[7] = a[0] ^ a[3] ^ a[6] ^ a[7];
            end
        8'd157:
            begin
                z[0] = a[0] ^ a[1] ^ a[4] ^ a[7];
                z[1] = a[1] ^ a[2] ^ a[5];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[5];
                z[4] = a[0] ^ a[3] ^ a[6] ^ a[7];
                z[5] = a[1] ^ a[4] ^ a[7];
                z[6] = a[2] ^ a[5];
                z[7] = a[0] ^ a[3] ^ a[6];
            end
        8'd158:
            begin
                z[0] = a[1] ^ a[4];
                z[1] = a[0] ^ a[2] ^ a[5];
                z[2] = a[0] ^ a[3] ^ a[4] ^ a[6];
                z[3] = a[0] ^ a[5] ^ a[7];
                z[4] = a[0] ^ a[4] ^ a[6];
                z[5] = a[1] ^ a[5] ^ a[7];
                z[6] = a[2] ^ a[6];
                z[7] = a[0] ^ a[3] ^ a[7];
            end
        8'd159:
            begin
                z[0] = a[0] ^ a[1] ^ a[4];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[5];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[3] = a[0] ^ a[3] ^ a[5] ^ a[7];
                z[4] = a[0] ^ a[6];
                z[5] = a[1] ^ a[7];
                z[6] = a[2];
                z[7] = a[0] ^ a[3];
            end
        8'd160:
            begin
                z[0] = a[1] ^ a[3] ^ a[5] ^ a[6];
                z[1] = a[2] ^ a[4] ^ a[6] ^ a[7];
                z[2] = a[1] ^ a[6] ^ a[7];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[5] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[6] = a[1] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
            end
        8'd161:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[6];
                z[1] = a[1] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[2] = a[1] ^ a[2] ^ a[6] ^ a[7];
                z[3] = a[1] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[1] ^ a[2] ^ a[5] ^ a[7];
                z[5] = a[0] ^ a[2] ^ a[3] ^ a[6];
                z[6] = a[1] ^ a[3] ^ a[4] ^ a[7];
                z[7] = a[0] ^ a[2] ^ a[4] ^ a[5];
            end
        8'd162:
            begin
                z[0] = a[1] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[2] = a[6];
                z[3] = a[1] ^ a[3] ^ a[5] ^ a[6];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[5] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd163:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[2] = a[2] ^ a[6];
                z[3] = a[1] ^ a[5] ^ a[6];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[5];
                z[5] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[6] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[7] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
            end
        8'd164:
            begin
                z[0] = a[1] ^ a[3] ^ a[5];
                z[1] = a[2] ^ a[4] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[7];
                z[3] = a[2] ^ a[3] ^ a[5];
                z[4] = a[1] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[1] ^ a[3] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[2] ^ a[4] ^ a[7];
            end
        8'd165:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[5];
                z[1] = a[1] ^ a[2] ^ a[4] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[7];
                z[3] = a[2] ^ a[5];
                z[4] = a[1] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[2] ^ a[6] ^ a[7];
                z[6] = a[1] ^ a[3] ^ a[7];
                z[7] = a[0] ^ a[2] ^ a[4];
            end
        8'd166:
            begin
                z[0] = a[1] ^ a[3] ^ a[5] ^ a[7];
                z[1] = a[0] ^ a[2] ^ a[4] ^ a[6];
                z[2] = a[0];
                z[3] = a[3] ^ a[5] ^ a[7];
                z[4] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[1] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
            end
        8'd167:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[6];
                z[2] = a[0] ^ a[2];
                z[3] = a[5] ^ a[7];
                z[4] = a[1] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[6] = a[1] ^ a[3] ^ a[5] ^ a[7];
                z[7] = a[0] ^ a[2] ^ a[4] ^ a[6];
            end
        8'd168:
            begin
                z[0] = a[1] ^ a[3] ^ a[6];
                z[1] = a[2] ^ a[4] ^ a[7];
                z[2] = a[1] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[7];
                z[4] = a[2] ^ a[4] ^ a[6];
                z[5] = a[0] ^ a[3] ^ a[5] ^ a[7];
                z[6] = a[1] ^ a[4] ^ a[6];
                z[7] = a[0] ^ a[2] ^ a[5] ^ a[7];
            end
        8'd169:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[6];
                z[1] = a[1] ^ a[2] ^ a[4] ^ a[7];
                z[2] = a[1] ^ a[2] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[7];
                z[4] = a[2] ^ a[6];
                z[5] = a[0] ^ a[3] ^ a[7];
                z[6] = a[1] ^ a[4];
                z[7] = a[0] ^ a[2] ^ a[5];
            end
        8'd170:
            begin
                z[0] = a[1] ^ a[3] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[2] ^ a[4] ^ a[7];
                z[2] = a[5] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[3];
                z[4] = a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[6] = a[1] ^ a[4] ^ a[5] ^ a[6];
                z[7] = a[0] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd171:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[7];
                z[2] = a[2] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[1];
                z[4] = a[2] ^ a[3] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[3] ^ a[4] ^ a[7];
                z[6] = a[1] ^ a[4] ^ a[5];
                z[7] = a[0] ^ a[2] ^ a[5] ^ a[6];
            end
        8'd172:
            begin
                z[0] = a[1] ^ a[3];
                z[1] = a[2] ^ a[4];
                z[2] = a[0] ^ a[1] ^ a[5];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[6];
                z[4] = a[4] ^ a[7];
                z[5] = a[0] ^ a[5];
                z[6] = a[1] ^ a[6];
                z[7] = a[0] ^ a[2] ^ a[7];
            end
        8'd173:
            begin
                z[0] = a[0] ^ a[1] ^ a[3];
                z[1] = a[1] ^ a[2] ^ a[4];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[5];
                z[3] = a[0] ^ a[2] ^ a[6];
                z[4] = a[7];
                z[5] = a[0];
                z[6] = a[1];
                z[7] = a[0] ^ a[2];
            end
        8'd174:
            begin
                z[0] = a[1] ^ a[3] ^ a[7];
                z[1] = a[0] ^ a[2] ^ a[4];
                z[2] = a[0] ^ a[5] ^ a[7];
                z[3] = a[0] ^ a[3] ^ a[6] ^ a[7];
                z[4] = a[3] ^ a[4];
                z[5] = a[0] ^ a[4] ^ a[5];
                z[6] = a[1] ^ a[5] ^ a[6];
                z[7] = a[0] ^ a[2] ^ a[6] ^ a[7];
            end
        8'd175:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[4];
                z[2] = a[0] ^ a[2] ^ a[5] ^ a[7];
                z[3] = a[0] ^ a[6] ^ a[7];
                z[4] = a[3];
                z[5] = a[0] ^ a[4];
                z[6] = a[1] ^ a[5];
                z[7] = a[0] ^ a[2] ^ a[6];
            end
        8'd176:
            begin
                z[0] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[1] ^ a[4] ^ a[7];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[7];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[4];
                z[7] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
            end
        8'd177:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[1] ^ a[2] ^ a[4] ^ a[7];
                z[3] = a[1] ^ a[2] ^ a[4] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[7] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
            end
        8'd178:
            begin
                z[0] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[4];
                z[3] = a[1] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[7] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
            end
        8'd179:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[2] ^ a[4];
                z[3] = a[1] ^ a[4] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[7] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd180:
            begin
                z[0] = a[1] ^ a[3] ^ a[4] ^ a[5];
                z[1] = a[2] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[4] ^ a[6] ^ a[7];
                z[3] = a[2] ^ a[3] ^ a[4] ^ a[7];
                z[4] = a[0] ^ a[1];
                z[5] = a[0] ^ a[1] ^ a[2];
                z[6] = a[1] ^ a[2] ^ a[3];
                z[7] = a[0] ^ a[2] ^ a[3] ^ a[4];
            end
        8'd181:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5];
                z[1] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[3] = a[2] ^ a[4] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[4];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[5];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[6];
                z[7] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
            end
        8'd182:
            begin
                z[0] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[1] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[4] ^ a[6];
                z[3] = a[3] ^ a[4];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[4];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[5];
                z[7] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
            end
        8'd183:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[0] ^ a[2] ^ a[4] ^ a[6];
                z[3] = a[4];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5];
                z[6] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[7] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
            end
        8'd184:
            begin
                z[0] = a[1] ^ a[3] ^ a[4] ^ a[6];
                z[1] = a[2] ^ a[4] ^ a[5] ^ a[7];
                z[2] = a[1] ^ a[4] ^ a[5];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[4] = a[0] ^ a[2] ^ a[5];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[6];
                z[6] = a[1] ^ a[2] ^ a[4] ^ a[7];
                z[7] = a[0] ^ a[2] ^ a[3] ^ a[5];
            end
        8'd185:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6];
                z[1] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[2] = a[1] ^ a[2] ^ a[4] ^ a[5];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5];
                z[4] = a[0] ^ a[2] ^ a[4] ^ a[5];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[6];
                z[6] = a[1] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
            end
        8'd186:
            begin
                z[0] = a[1] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[2] = a[4] ^ a[5] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6];
                z[6] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[7] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
            end
        8'd187:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[2] = a[2] ^ a[4] ^ a[5] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[7];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd188:
            begin
                z[0] = a[1] ^ a[3] ^ a[4];
                z[1] = a[2] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[6] ^ a[7];
                z[6] = a[1] ^ a[2] ^ a[7];
                z[7] = a[0] ^ a[2] ^ a[3];
            end
        8'd189:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[4];
                z[1] = a[1] ^ a[2] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[1] ^ a[2] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[2] ^ a[3] ^ a[7];
            end
        8'd190:
            begin
                z[0] = a[1] ^ a[3] ^ a[4] ^ a[7];
                z[1] = a[0] ^ a[2] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[3] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[4] ^ a[6] ^ a[7];
                z[6] = a[1] ^ a[2] ^ a[5] ^ a[7];
                z[7] = a[0] ^ a[2] ^ a[3] ^ a[6];
            end
        8'd191:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5];
                z[2] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[1] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
            end
        8'd192:
            begin
                z[0] = a[1] ^ a[2] ^ a[5];
                z[1] = a[2] ^ a[3] ^ a[6];
                z[2] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[3] = a[1] ^ a[3] ^ a[4] ^ a[6];
                z[4] = a[1] ^ a[4] ^ a[7];
                z[5] = a[2] ^ a[5];
                z[6] = a[0] ^ a[3] ^ a[6];
                z[7] = a[0] ^ a[1] ^ a[4] ^ a[7];
            end
        8'd193:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[5];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[6];
                z[2] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[3] = a[1] ^ a[4] ^ a[6];
                z[4] = a[1] ^ a[7];
                z[5] = a[2];
                z[6] = a[0] ^ a[3];
                z[7] = a[0] ^ a[1] ^ a[4];
            end
        8'd194:
            begin
                z[0] = a[1] ^ a[2] ^ a[5] ^ a[7];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[6];
                z[2] = a[2] ^ a[3] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[4] = a[1] ^ a[3] ^ a[4];
                z[5] = a[2] ^ a[4] ^ a[5];
                z[6] = a[0] ^ a[3] ^ a[5] ^ a[6];
                z[7] = a[0] ^ a[1] ^ a[4] ^ a[6] ^ a[7];
            end
        8'd195:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6];
                z[2] = a[3] ^ a[4] ^ a[5];
                z[3] = a[1] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[4] = a[1] ^ a[3];
                z[5] = a[2] ^ a[4];
                z[6] = a[0] ^ a[3] ^ a[5];
                z[7] = a[0] ^ a[1] ^ a[4] ^ a[6];
            end
        8'd196:
            begin
                z[0] = a[1] ^ a[2] ^ a[5] ^ a[6];
                z[1] = a[2] ^ a[3] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[3] ^ a[4] ^ a[7];
                z[4] = a[1] ^ a[2] ^ a[4] ^ a[6];
                z[5] = a[2] ^ a[3] ^ a[5] ^ a[7];
                z[6] = a[0] ^ a[3] ^ a[4] ^ a[6];
                z[7] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[7];
            end
        8'd197:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[4] ^ a[7];
                z[4] = a[1] ^ a[2] ^ a[6];
                z[5] = a[2] ^ a[3] ^ a[7];
                z[6] = a[0] ^ a[3] ^ a[4];
                z[7] = a[0] ^ a[1] ^ a[4] ^ a[5];
            end
        8'd198:
            begin
                z[0] = a[1] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[2] ^ a[3] ^ a[4];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[5] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[6] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[7] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd199:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[2] ^ a[4];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[5] = a[2] ^ a[3] ^ a[4] ^ a[7];
                z[6] = a[0] ^ a[3] ^ a[4] ^ a[5];
                z[7] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6];
            end
        8'd200:
            begin
                z[0] = a[1] ^ a[2];
                z[1] = a[2] ^ a[3];
                z[2] = a[1] ^ a[2] ^ a[3] ^ a[4];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5];
                z[4] = a[4] ^ a[5] ^ a[6];
                z[5] = a[5] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[7];
            end
        8'd201:
            begin
                z[0] = a[0] ^ a[1] ^ a[2];
                z[1] = a[1] ^ a[2] ^ a[3];
                z[2] = a[1] ^ a[3] ^ a[4];
                z[3] = a[0] ^ a[1] ^ a[4] ^ a[5];
                z[4] = a[5] ^ a[6];
                z[5] = a[6] ^ a[7];
                z[6] = a[0] ^ a[7];
                z[7] = a[0] ^ a[1];
            end
        8'd202:
            begin
                z[0] = a[1] ^ a[2] ^ a[7];
                z[1] = a[0] ^ a[2] ^ a[3];
                z[2] = a[2] ^ a[3] ^ a[4] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[4] = a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[4] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[6] ^ a[7];
            end
        8'd203:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3];
                z[2] = a[3] ^ a[4] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[4] = a[3] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[4] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[5] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[6];
            end
        8'd204:
            begin
                z[0] = a[1] ^ a[2] ^ a[6];
                z[1] = a[2] ^ a[3] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[3] = a[0] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[2] ^ a[4] ^ a[5] ^ a[7];
                z[5] = a[3] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[4] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[5] ^ a[7];
            end
        8'd205:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[6];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6];
                z[3] = a[0] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[2] ^ a[5] ^ a[7];
                z[5] = a[3] ^ a[6];
                z[6] = a[0] ^ a[4] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[5];
            end
        8'd206:
            begin
                z[0] = a[1] ^ a[2] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[7];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[2] ^ a[3] ^ a[4] ^ a[5];
                z[5] = a[3] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd207:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[7];
                z[2] = a[0] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[2] ^ a[3] ^ a[5];
                z[5] = a[3] ^ a[4] ^ a[6];
                z[6] = a[0] ^ a[4] ^ a[5] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[5] ^ a[6];
            end
        8'd208:
            begin
                z[0] = a[1] ^ a[2] ^ a[4] ^ a[5];
                z[1] = a[2] ^ a[3] ^ a[5] ^ a[6];
                z[2] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[1] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[1] ^ a[2] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[2] ^ a[3] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[3] ^ a[4];
            end
        8'd209:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[2] = a[1] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[1] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[1] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[7];
            end
        8'd210:
            begin
                z[0] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[2] = a[2] ^ a[3] ^ a[5] ^ a[6];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[6];
                z[5] = a[1] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6];
            end
        8'd211:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[2] = a[3] ^ a[5] ^ a[6];
                z[3] = a[1] ^ a[2] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
            end
        8'd212:
            begin
                z[0] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[3] = a[3] ^ a[5];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[5];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[6];
                z[6] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5];
            end
        8'd213:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[7];
                z[3] = a[5];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
            end
        8'd214:
            begin
                z[0] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[5];
                z[3] = a[2] ^ a[3] ^ a[5] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[6] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
            end
        8'd215:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[3] ^ a[5];
                z[3] = a[2] ^ a[5] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[5] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd216:
            begin
                z[0] = a[1] ^ a[2] ^ a[4];
                z[1] = a[2] ^ a[3] ^ a[5];
                z[2] = a[1] ^ a[2] ^ a[3] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[7];
                z[4] = a[0];
                z[5] = a[1];
                z[6] = a[0] ^ a[2];
                z[7] = a[0] ^ a[1] ^ a[3];
            end
        8'd217:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[4];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[5];
                z[2] = a[1] ^ a[3] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[7];
                z[4] = a[0] ^ a[4];
                z[5] = a[1] ^ a[5];
                z[6] = a[0] ^ a[2] ^ a[6];
                z[7] = a[0] ^ a[1] ^ a[3] ^ a[7];
            end
        8'd218:
            begin
                z[0] = a[1] ^ a[2] ^ a[4] ^ a[7];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[5];
                z[2] = a[2] ^ a[3] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3];
                z[4] = a[0] ^ a[3] ^ a[7];
                z[5] = a[1] ^ a[4];
                z[6] = a[0] ^ a[2] ^ a[5];
                z[7] = a[0] ^ a[1] ^ a[3] ^ a[6];
            end
        8'd219:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5];
                z[2] = a[3] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[2];
                z[4] = a[0] ^ a[3] ^ a[4] ^ a[7];
                z[5] = a[1] ^ a[4] ^ a[5];
                z[6] = a[0] ^ a[2] ^ a[5] ^ a[6];
                z[7] = a[0] ^ a[1] ^ a[3] ^ a[6] ^ a[7];
            end
        8'd220:
            begin
                z[0] = a[1] ^ a[2] ^ a[4] ^ a[6];
                z[1] = a[2] ^ a[3] ^ a[5] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3];
                z[3] = a[0] ^ a[3] ^ a[6];
                z[4] = a[0] ^ a[2] ^ a[6] ^ a[7];
                z[5] = a[1] ^ a[3] ^ a[7];
                z[6] = a[0] ^ a[2] ^ a[4];
                z[7] = a[0] ^ a[1] ^ a[3] ^ a[5];
            end
        8'd221:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[6];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[3];
                z[3] = a[0] ^ a[6];
                z[4] = a[0] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[5] = a[1] ^ a[3] ^ a[5] ^ a[7];
                z[6] = a[0] ^ a[2] ^ a[4] ^ a[6];
                z[7] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[7];
            end
        8'd222:
            begin
                z[0] = a[1] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[2] = a[0] ^ a[2] ^ a[3] ^ a[7];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[6];
                z[5] = a[1] ^ a[3] ^ a[4] ^ a[7];
                z[6] = a[0] ^ a[2] ^ a[4] ^ a[5];
                z[7] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[6];
            end
        8'd223:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[2] = a[0] ^ a[3] ^ a[7];
                z[3] = a[0] ^ a[2] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[5] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[6] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[7] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd224:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[1] = a[2] ^ a[3] ^ a[4] ^ a[6];
                z[2] = a[1] ^ a[2] ^ a[4];
                z[3] = a[1] ^ a[7];
                z[4] = a[1] ^ a[3] ^ a[5] ^ a[7];
                z[5] = a[0] ^ a[2] ^ a[4] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[6];
            end
        8'd225:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[2] = a[1] ^ a[4];
                z[3] = a[1] ^ a[3] ^ a[7];
                z[4] = a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[5] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
            end
        8'd226:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[5];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[2] = a[2] ^ a[4] ^ a[7];
                z[3] = a[1] ^ a[2];
                z[4] = a[1] ^ a[5];
                z[5] = a[0] ^ a[2] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[3] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[4];
            end
        8'd227:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[2] = a[4] ^ a[7];
                z[3] = a[1] ^ a[2] ^ a[3];
                z[4] = a[1] ^ a[4] ^ a[5];
                z[5] = a[0] ^ a[2] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[3] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[7];
            end
        8'd228:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[6];
                z[3] = a[6];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
            end
        8'd229:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[4] ^ a[6];
                z[3] = a[3] ^ a[6];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd230:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[3] = a[2] ^ a[6] ^ a[7];
                z[4] = a[1] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5];
            end
        8'd231:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[4] ^ a[6] ^ a[7];
                z[3] = a[2] ^ a[3] ^ a[6] ^ a[7];
                z[4] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
            end
        8'd232:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[7];
                z[1] = a[2] ^ a[3] ^ a[4];
                z[2] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[3] ^ a[6];
                z[5] = a[0] ^ a[4] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[5];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[6];
            end
        8'd233:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[7];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[4];
                z[2] = a[1] ^ a[4] ^ a[5] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[3] ^ a[4] ^ a[6];
                z[5] = a[0] ^ a[4] ^ a[5] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[5] ^ a[6];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[6] ^ a[7];
            end
        8'd234:
            begin
                z[0] = a[1] ^ a[2] ^ a[3];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[2] = a[2] ^ a[4] ^ a[5];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6];
                z[4] = a[6] ^ a[7];
                z[5] = a[0] ^ a[7];
                z[6] = a[0] ^ a[1];
                z[7] = a[0] ^ a[1] ^ a[2];
            end
        8'd235:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
                z[2] = a[4] ^ a[5];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[4] = a[4] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[5] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[6];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[7];
            end
        8'd236:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[1] = a[2] ^ a[3] ^ a[4] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[5];
                z[4] = a[2] ^ a[3] ^ a[7];
                z[5] = a[0] ^ a[3] ^ a[4];
                z[6] = a[0] ^ a[1] ^ a[4] ^ a[5];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6];
            end
        8'd237:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[3] ^ a[5];
                z[4] = a[2] ^ a[3] ^ a[4] ^ a[7];
                z[5] = a[0] ^ a[3] ^ a[4] ^ a[5];
                z[6] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd238:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[6];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[2] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[2] ^ a[5] ^ a[7];
                z[4] = a[2];
                z[5] = a[0] ^ a[3];
                z[6] = a[0] ^ a[1] ^ a[4];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[5];
            end
        8'd239:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[2] = a[0] ^ a[4] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
                z[4] = a[2] ^ a[4];
                z[5] = a[0] ^ a[3] ^ a[5];
                z[6] = a[0] ^ a[1] ^ a[4] ^ a[6];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[7];
            end
        8'd240:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[1] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[1] ^ a[2] ^ a[6];
                z[3] = a[1] ^ a[4] ^ a[5];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
            end
        8'd241:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[1] ^ a[6];
                z[3] = a[1] ^ a[3] ^ a[4] ^ a[5];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
            end
        8'd242:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[2] ^ a[6] ^ a[7];
                z[3] = a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[4] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
            end
        8'd243:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[2] = a[6] ^ a[7];
                z[3] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
            end
        8'd244:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[2];
                z[3] = a[4] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd245:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[1];
                z[3] = a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
            end
        8'd246:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[2] ^ a[7];
                z[3] = a[2] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
            end
        8'd247:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[2] = a[0] ^ a[7];
                z[3] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[2] ^ a[3];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
            end
        8'd248:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[1] = a[2] ^ a[3] ^ a[4] ^ a[5];
                z[2] = a[1] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[4] ^ a[6];
                z[4] = a[0] ^ a[3] ^ a[4] ^ a[5];
                z[5] = a[0] ^ a[1] ^ a[4] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6] ^ a[7];
            end
        8'd249:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[7];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[2] = a[1] ^ a[5] ^ a[6] ^ a[7];
                z[3] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6];
                z[4] = a[0] ^ a[3] ^ a[5];
                z[5] = a[0] ^ a[1] ^ a[4] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[6];
            end
        8'd250:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[4];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[2] = a[2] ^ a[5] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[4] ^ a[5] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[5] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[7];
            end
        8'd251:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5];
                z[2] = a[5] ^ a[6];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[4] = a[0] ^ a[5] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[6];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[3];
            end
        8'd252:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[1] = a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[5] ^ a[7];
                z[3] = a[0] ^ a[4] ^ a[7];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
            end
        8'd253:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[2] = a[0] ^ a[1] ^ a[5] ^ a[7];
                z[3] = a[0] ^ a[3] ^ a[4] ^ a[7];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[4] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[5] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[6];
            end
        8'd254:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[2] = a[0] ^ a[2] ^ a[5];
                z[3] = a[0] ^ a[2] ^ a[4];
                z[4] = a[0] ^ a[2] ^ a[4] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[5] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[6] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5] ^ a[7];
            end
        8'd255:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[6];
                z[1] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4] ^ a[5] ^ a[7];
                z[2] = a[0] ^ a[5];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[4] = a[0] ^ a[2] ^ a[5] ^ a[6];
                z[5] = a[0] ^ a[1] ^ a[3] ^ a[6] ^ a[7];
                z[6] = a[0] ^ a[1] ^ a[2] ^ a[4] ^ a[7];
                z[7] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[5];
            end
        default:
            begin
                z[0] = 0; 
                z[1] = 0; 
                z[2] = 0; 
                z[3] = 0; 
                z[4] = 0; 
                z[5] = 0; 
                z[6] = 0; 
                z[7] = 0; 
            end
    endcase
end
endmodule
