//`include "hpilot_preprocess_if.sv"  

`include "smp_if.sv" 
`include "test_collection_enc.sv" 