
`timescale 1ns/100ps

module kes #( parameter [
`SYM_BW_BW -1 :0] SYM_BW = 8,

parameter [8-1:0]  N_NUM = 255, parameter [
`R_BW - 1 :0]  R_NUM = 16,

parameter [
`R_BW - 1 :0]  T_NUM = R_NUM/2

)  (        input clk,        input rst_n,        input start,         input [SYM_BW*R_NUM - 1:0] syndrome   ,        output reg [SYM_BW*(T_NUM+1) - 1:0] lamda,        output reg [SYM_BW*(T_NUM) - 1:0] omega,                  output reg done         );     reg [SYM_BW-1:0] ID_S_f49cf8f_3369e3c5_E[3*T_NUM+1:0]; reg [SYM_BW-1:0] ID_S_106cdefb_6c58346a_E[3*T_NUM  :0]; reg signed [7:0] ID_S_7c995d3e_78e7367b_E        ; reg [SYM_BW-1:0] ID_S_f7deae8_3b9c8f15_E       ; reg [7:0] ID_S_651d5efd_799ab730_E       ;  reg ID_S_354d19ab_1a25e150_E;    wire [SYM_BW-1:0] ID_S_16c253ca_7bef0f84_E[3*T_NUM  :0]; wire [SYM_BW-1:0] ID_S_1949e91d_47b560eb_E[3*T_NUM  :0];   always @(posedge clk or negedge rst_n) if (!rst_n)   ID_S_651d5efd_799ab730_E <= 8'd0; else if (start)   ID_S_651d5efd_799ab730_E <= 8'd1; else if ((ID_S_651d5efd_799ab730_E < 2*T_NUM ) && ID_S_651d5efd_799ab730_E)   ID_S_651d5efd_799ab730_E <= ID_S_651d5efd_799ab730_E + 8'd1; else    ID_S_651d5efd_799ab730_E <= 8'd0;     always @(posedge clk or negedge rst_n) if (!rst_n)   ID_S_354d19ab_1a25e150_E <= 1'd0; else if (ID_S_651d5efd_799ab730_E == 2*T_NUM)   ID_S_354d19ab_1a25e150_E <= 1'd1; else    ID_S_354d19ab_1a25e150_E <= 1'd0;    genvar ID_S_37eae313_2f21b4b4_E; generate     for(ID_S_37eae313_2f21b4b4_E = 0;ID_S_37eae313_2f21b4b4_E <= 2*T_NUM - 1 ;ID_S_37eae313_2f21b4b4_E = ID_S_37eae313_2f21b4b4_E + 1)     begin         always @(posedge clk or negedge rst_n)         if (!rst_n)             begin                 ID_S_f49cf8f_3369e3c5_E[ID_S_37eae313_2f21b4b4_E]       <= {SYM_BW{1'b0}};               end         else if (start)             begin                 ID_S_f49cf8f_3369e3c5_E[ID_S_37eae313_2f21b4b4_E]       <= syndrome[(ID_S_37eae313_2f21b4b4_E+1) *SYM_BW - 1:ID_S_37eae313_2f21b4b4_E *SYM_BW] ;               end             else if(ID_S_651d5efd_799ab730_E)             begin                 ID_S_f49cf8f_3369e3c5_E[ID_S_37eae313_2f21b4b4_E]       <= ID_S_16c253ca_7bef0f84_E[ID_S_37eae313_2f21b4b4_E]       ^ ID_S_1949e91d_47b560eb_E[ID_S_37eae313_2f21b4b4_E]   ;              end         else             begin                 ID_S_f49cf8f_3369e3c5_E[ID_S_37eae313_2f21b4b4_E]       <= {SYM_BW{1'b0}};               end             end endgenerate  generate     for(ID_S_37eae313_2f21b4b4_E = 2*T_NUM ;ID_S_37eae313_2f21b4b4_E <= 3*T_NUM - 1 ;ID_S_37eae313_2f21b4b4_E = ID_S_37eae313_2f21b4b4_E + 1)     begin         always @(posedge clk or negedge rst_n)         if (!rst_n)             begin                 ID_S_f49cf8f_3369e3c5_E[ID_S_37eae313_2f21b4b4_E]       <= {SYM_BW{1'b0}};               end         else if (start)             begin                 ID_S_f49cf8f_3369e3c5_E[ID_S_37eae313_2f21b4b4_E]       <= {SYM_BW{1'b0}};             end         else if(ID_S_651d5efd_799ab730_E)             begin                             ID_S_f49cf8f_3369e3c5_E[ID_S_37eae313_2f21b4b4_E]       <= ID_S_16c253ca_7bef0f84_E[ID_S_37eae313_2f21b4b4_E]       ^ ID_S_1949e91d_47b560eb_E[ID_S_37eae313_2f21b4b4_E]   ;              end         else             begin                 ID_S_f49cf8f_3369e3c5_E[ID_S_37eae313_2f21b4b4_E]       <= {SYM_BW{1'b0}};               end             end endgenerate  always @(posedge clk or negedge rst_n) if (!rst_n)     ID_S_f49cf8f_3369e3c5_E[3*T_NUM]       <= {SYM_BW{1'b0}}; else if (start)         ID_S_f49cf8f_3369e3c5_E[3*T_NUM]       <= {{(SYM_BW-1){1'b0}},{1'b1}}; else if(ID_S_651d5efd_799ab730_E)     ID_S_f49cf8f_3369e3c5_E[3*T_NUM]       <= ID_S_16c253ca_7bef0f84_E[3*T_NUM]       ^ ID_S_1949e91d_47b560eb_E[3*T_NUM]   ;  else     ID_S_f49cf8f_3369e3c5_E[3*T_NUM] <= 0;    always @(posedge clk or negedge rst_n) if (!rst_n)         ID_S_f49cf8f_3369e3c5_E[3*T_NUM+1]       <= {SYM_BW{1'b0}}; else if (start)         ID_S_f49cf8f_3369e3c5_E[3*T_NUM+1]       <= {SYM_BW{1'b0}}; else ;   genvar ID_S_299fc87f_25d392ef_E; generate     for(ID_S_299fc87f_25d392ef_E = 0;ID_S_299fc87f_25d392ef_E <= 2*T_NUM - 1 ;ID_S_299fc87f_25d392ef_E = ID_S_299fc87f_25d392ef_E + 1)     begin         always @(posedge clk or negedge rst_n)         if (!rst_n)             begin                 ID_S_106cdefb_6c58346a_E[ID_S_299fc87f_25d392ef_E]       <= {SYM_BW{1'b0}};               end         else if (start)             begin                 ID_S_106cdefb_6c58346a_E[ID_S_299fc87f_25d392ef_E]       <= syndrome[(ID_S_299fc87f_25d392ef_E+1) *SYM_BW - 1:ID_S_299fc87f_25d392ef_E *SYM_BW] ;               end             else if(ID_S_651d5efd_799ab730_E)         begin           if((ID_S_f49cf8f_3369e3c5_E[0]) && (ID_S_7c995d3e_78e7367b_E >= 0)) begin               ID_S_106cdefb_6c58346a_E[ID_S_299fc87f_25d392ef_E]         <= ID_S_f49cf8f_3369e3c5_E[ID_S_299fc87f_25d392ef_E+1      ];           end else             ;          end         else             begin                 ID_S_106cdefb_6c58346a_E[ID_S_299fc87f_25d392ef_E]       <= {SYM_BW{1'b0}};             end     end endgenerate  generate     for(ID_S_299fc87f_25d392ef_E = 2*T_NUM;ID_S_299fc87f_25d392ef_E <= 3*T_NUM - 1 ;ID_S_299fc87f_25d392ef_E = ID_S_299fc87f_25d392ef_E + 1)     begin         always @(posedge clk or negedge rst_n)         if (!rst_n)             begin                 ID_S_106cdefb_6c58346a_E[ID_S_299fc87f_25d392ef_E]       <= {SYM_BW{1'b0}};              end         else if (start)             begin                 ID_S_106cdefb_6c58346a_E[ID_S_299fc87f_25d392ef_E]       <= {SYM_BW{1'b0}};             end             else if(ID_S_651d5efd_799ab730_E)         begin           if((ID_S_f49cf8f_3369e3c5_E[0]) && (ID_S_7c995d3e_78e7367b_E >= 0)) begin               ID_S_106cdefb_6c58346a_E[ID_S_299fc87f_25d392ef_E      ]     <= ID_S_f49cf8f_3369e3c5_E[ID_S_299fc87f_25d392ef_E+1      ];           end else             ;          end         else             begin                 ID_S_106cdefb_6c58346a_E[ID_S_299fc87f_25d392ef_E]       <= {SYM_BW{1'b0}};              end             end endgenerate  always @(posedge clk or negedge rst_n) if (!rst_n)     begin         ID_S_106cdefb_6c58346a_E[3*T_NUM]       <= {SYM_BW{1'b0}};     end else if (start)     begin         ID_S_106cdefb_6c58346a_E[3*T_NUM]       <= {{(SYM_BW-1){1'b0}},{1'b1}};     end     else if(ID_S_651d5efd_799ab730_E)     begin       if((ID_S_f49cf8f_3369e3c5_E[0]) && (ID_S_7c995d3e_78e7367b_E >= 0)) begin           ID_S_106cdefb_6c58346a_E[3*T_NUM      ]     <= ID_S_f49cf8f_3369e3c5_E[3*T_NUM+1      ];       end else         ;      end  else     ID_S_106cdefb_6c58346a_E[3*T_NUM]       <= {SYM_BW{1'b0}};    always @(posedge clk or negedge rst_n) if (!rst_n)     begin         ID_S_7c995d3e_78e7367b_E  <= 8'd0;         ID_S_f7deae8_3b9c8f15_E <= {SYM_BW{1'b0}};     end else if(start)     begin         ID_S_7c995d3e_78e7367b_E  <= 8'd0;         ID_S_f7deae8_3b9c8f15_E <= {{(SYM_BW-1){1'b0}},{1'b1}};     end else if(ID_S_651d5efd_799ab730_E )     begin         if((ID_S_f49cf8f_3369e3c5_E[0] ) && (ID_S_7c995d3e_78e7367b_E >= 0)) begin             ID_S_f7deae8_3b9c8f15_E <= ID_S_f49cf8f_3369e3c5_E[0];             ID_S_7c995d3e_78e7367b_E  <= -ID_S_7c995d3e_78e7367b_E - 1;         end else begin             ID_S_f7deae8_3b9c8f15_E <= ID_S_f7deae8_3b9c8f15_E;             ID_S_7c995d3e_78e7367b_E  <= ID_S_7c995d3e_78e7367b_E+1;         end     end else     begin         ID_S_7c995d3e_78e7367b_E  <= 8'd0;         ID_S_f7deae8_3b9c8f15_E <= {{(SYM_BW-1){1'b0}},{1'b1}};     end  generate     for(ID_S_299fc87f_25d392ef_E = 0;ID_S_299fc87f_25d392ef_E <= 3*T_NUM  ;ID_S_299fc87f_25d392ef_E = ID_S_299fc87f_25d392ef_E + 1)     begin         case({SYM_BW})             {4'd3}:             begin:gf8mul_dec                 gf8mul_dec   ID_S_60071ffb_49a40e8d_E( ID_S_f49cf8f_3369e3c5_E[ID_S_299fc87f_25d392ef_E+1] ,  ID_S_f7deae8_3b9c8f15_E            ,  ID_S_16c253ca_7bef0f84_E[ID_S_299fc87f_25d392ef_E] );                 gf8mul_dec   ID_S_6019387c_49564b10_E( ID_S_f49cf8f_3369e3c5_E[0]           ,  ID_S_106cdefb_6c58346a_E[ID_S_299fc87f_25d392ef_E] ,  ID_S_1949e91d_47b560eb_E[ID_S_299fc87f_25d392ef_E] );                        end                                                                                                                                                                                                                 {4'd4}:                                                                                                   begin:gf16mul_dec                                                                                             gf16mul_dec  ID_S_60071ffb_49a40e8d_E( ID_S_f49cf8f_3369e3c5_E[ID_S_299fc87f_25d392ef_E+1] ,  ID_S_f7deae8_3b9c8f15_E            ,  ID_S_16c253ca_7bef0f84_E[ID_S_299fc87f_25d392ef_E] );                 gf16mul_dec  ID_S_6019387c_49564b10_E( ID_S_f49cf8f_3369e3c5_E[0]           ,  ID_S_106cdefb_6c58346a_E[ID_S_299fc87f_25d392ef_E] ,  ID_S_1949e91d_47b560eb_E[ID_S_299fc87f_25d392ef_E] );                        end                                                                                                                                                                                                                 {4'd5}:                                                                                                   begin:gf32mul_dec                                                                                             gf32mul_dec  ID_S_60071ffb_49a40e8d_E( ID_S_f49cf8f_3369e3c5_E[ID_S_299fc87f_25d392ef_E+1] ,  ID_S_f7deae8_3b9c8f15_E            ,  ID_S_16c253ca_7bef0f84_E[ID_S_299fc87f_25d392ef_E] );                 gf32mul_dec  ID_S_6019387c_49564b10_E( ID_S_f49cf8f_3369e3c5_E[0]           ,  ID_S_106cdefb_6c58346a_E[ID_S_299fc87f_25d392ef_E] ,  ID_S_1949e91d_47b560eb_E[ID_S_299fc87f_25d392ef_E] );                        end                                                                                                                                                                                                                 {4'd6}:                                                                                                   begin:gf64mul_dec                                                                                             gf64mul_dec  ID_S_60071ffb_49a40e8d_E( ID_S_f49cf8f_3369e3c5_E[ID_S_299fc87f_25d392ef_E+1] ,  ID_S_f7deae8_3b9c8f15_E            ,  ID_S_16c253ca_7bef0f84_E[ID_S_299fc87f_25d392ef_E] );                 gf64mul_dec  ID_S_6019387c_49564b10_E( ID_S_f49cf8f_3369e3c5_E[0]           ,  ID_S_106cdefb_6c58346a_E[ID_S_299fc87f_25d392ef_E] ,  ID_S_1949e91d_47b560eb_E[ID_S_299fc87f_25d392ef_E] );                        end                                                                                                                                                                                                                 {4'd7}:                                                                                                   begin:gf128mul_dec                                                                                            gf128mul_dec ID_S_60071ffb_49a40e8d_E( ID_S_f49cf8f_3369e3c5_E[ID_S_299fc87f_25d392ef_E+1] ,  ID_S_f7deae8_3b9c8f15_E            ,  ID_S_16c253ca_7bef0f84_E[ID_S_299fc87f_25d392ef_E] );                 gf128mul_dec ID_S_6019387c_49564b10_E( ID_S_f49cf8f_3369e3c5_E[0]           ,  ID_S_106cdefb_6c58346a_E[ID_S_299fc87f_25d392ef_E] ,  ID_S_1949e91d_47b560eb_E[ID_S_299fc87f_25d392ef_E] );                        end                                                                                                                                                                                                                                                                                                                           {4'd8}:                                                                                                   begin:gf256mul_dec                                                                                            gf256mul_dec ID_S_60071ffb_49a40e8d_E( ID_S_f49cf8f_3369e3c5_E[ID_S_299fc87f_25d392ef_E+1] ,  ID_S_f7deae8_3b9c8f15_E            ,  ID_S_16c253ca_7bef0f84_E[ID_S_299fc87f_25d392ef_E] );                 gf256mul_dec ID_S_6019387c_49564b10_E( ID_S_f49cf8f_3369e3c5_E[0]           ,  ID_S_106cdefb_6c58346a_E[ID_S_299fc87f_25d392ef_E] ,  ID_S_1949e91d_47b560eb_E[ID_S_299fc87f_25d392ef_E] );             end         endcase                    end endgenerate    genvar ID_S_526eca48_36158cfe_E; generate     for(ID_S_526eca48_36158cfe_E = 0;ID_S_526eca48_36158cfe_E <= T_NUM  ;ID_S_526eca48_36158cfe_E = ID_S_526eca48_36158cfe_E + 1)     begin         always @(posedge clk or negedge rst_n)         if (!rst_n) begin                 lamda[(ID_S_526eca48_36158cfe_E+1) *SYM_BW - 1:ID_S_526eca48_36158cfe_E *SYM_BW]  <= 0;           end else if (ID_S_354d19ab_1a25e150_E) begin                         lamda[(ID_S_526eca48_36158cfe_E+1) *SYM_BW - 1:ID_S_526eca48_36158cfe_E *SYM_BW]   <= ID_S_f49cf8f_3369e3c5_E[T_NUM + ID_S_526eca48_36158cfe_E];                       end else ;     end endgenerate    genvar ID_S_6227abb2_151191de_E; generate     for(ID_S_6227abb2_151191de_E = 0;ID_S_6227abb2_151191de_E < T_NUM  ;ID_S_6227abb2_151191de_E = ID_S_6227abb2_151191de_E + 1)     begin         always @(posedge clk or negedge rst_n)         if (!rst_n) begin             omega[(ID_S_6227abb2_151191de_E + 1) *SYM_BW - 1:ID_S_6227abb2_151191de_E *SYM_BW]  <= 0;           end else if (ID_S_354d19ab_1a25e150_E) begin           omega[(ID_S_6227abb2_151191de_E + 1) *SYM_BW - 1:ID_S_6227abb2_151191de_E *SYM_BW]  <= ID_S_f49cf8f_3369e3c5_E[ ID_S_6227abb2_151191de_E];           end else            ;     end endgenerate     always @(posedge clk or negedge rst_n) if (!rst_n)     done  <= 1'b0; else     done  <= ID_S_354d19ab_1a25e150_E;   endmodule