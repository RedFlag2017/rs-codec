
`timescale 1ns/100ps

module err_locate #( parameter [
`SYM_BW_BW -1 :0] SYM_BW = 8,

parameter [8-1:0]  N_NUM = 255, parameter [
`R_BW - 1 :0]  R_NUM = 16,

parameter [
`R_BW - 1 :0]  T_NUM = R_NUM/2

)  (        input clk,        input rst_n,        input start,                 input [SYM_BW*(T_NUM+1) - 1:0] lamda,             output reg [SYM_BW*T_NUM - 1:0] err_loc    ,               output reg done        );          localparam [8 - 1 :0]  ID_S_53b735b7_11413ceb_E = 2**SYM_BW-1-N_NUM;        reg ID_S_787e79a3_1d07dd47_E; reg [4:0] ID_S_6f264d33_7f0e6051_E; reg [7:0] ID_S_651d5efd_799ab730_E;   wire [SYM_BW-1:0] ID_S_32a32f8d_795a5f17_E[2**SYM_BW-2:0]  ;  generate     case({SYM_BW})           4'd3:            begin               assign ID_S_32a32f8d_795a5f17_E[ 0]  = 3'd2;                assign ID_S_32a32f8d_795a5f17_E[ 1]  = 3'd4;                assign ID_S_32a32f8d_795a5f17_E[ 2]  = 3'd3;              assign ID_S_32a32f8d_795a5f17_E[ 3]  = 3'd6;              assign ID_S_32a32f8d_795a5f17_E[ 4]  = 3'd7;              assign ID_S_32a32f8d_795a5f17_E[ 5]  = 3'd5;              assign ID_S_32a32f8d_795a5f17_E[ 6]  = 3'd1;                            end         4'd4:            begin                  assign ID_S_32a32f8d_795a5f17_E[0 ]  =  4'd2;                 assign ID_S_32a32f8d_795a5f17_E[1 ]  =  4'd4;                 assign ID_S_32a32f8d_795a5f17_E[2 ]  =  4'd8;                 assign ID_S_32a32f8d_795a5f17_E[3 ]  =  4'd3;                  assign ID_S_32a32f8d_795a5f17_E[4 ]  =  4'd6;                 assign ID_S_32a32f8d_795a5f17_E[5 ]  =  4'd12;                 assign ID_S_32a32f8d_795a5f17_E[6 ]  =  4'd11;                 assign ID_S_32a32f8d_795a5f17_E[7 ]  =  4'd5;                 assign ID_S_32a32f8d_795a5f17_E[8 ]  =  4'd10;                 assign ID_S_32a32f8d_795a5f17_E[9 ]  =  4'd7;                 assign ID_S_32a32f8d_795a5f17_E[10]  =  4'd14;                 assign ID_S_32a32f8d_795a5f17_E[11]  =  4'd15;                 assign ID_S_32a32f8d_795a5f17_E[12]  =  4'd13;                 assign ID_S_32a32f8d_795a5f17_E[13]  =  4'd9;                 assign ID_S_32a32f8d_795a5f17_E[14]  =  4'd1;                       end         4'd5:            begin                  assign ID_S_32a32f8d_795a5f17_E[  0]  =  5'd2;                 assign ID_S_32a32f8d_795a5f17_E[  1]  =  5'd4;                 assign ID_S_32a32f8d_795a5f17_E[  2]  =  5'd8;                 assign ID_S_32a32f8d_795a5f17_E[  3]  =  5'd16;                  assign ID_S_32a32f8d_795a5f17_E[  4]  =  5'd5;                 assign ID_S_32a32f8d_795a5f17_E[  5]  =  5'd10;                 assign ID_S_32a32f8d_795a5f17_E[  6]  =  5'd20;                 assign ID_S_32a32f8d_795a5f17_E[  7]  =  5'd13;                  assign ID_S_32a32f8d_795a5f17_E[  8]  =  5'd26;                 assign ID_S_32a32f8d_795a5f17_E[  9]  =  5'd17;                 assign ID_S_32a32f8d_795a5f17_E[ 10]  =  5'd7;                 assign ID_S_32a32f8d_795a5f17_E[ 11]  =  5'd14;                  assign ID_S_32a32f8d_795a5f17_E[ 12]  =  5'd28;                 assign ID_S_32a32f8d_795a5f17_E[ 13]  =  5'd29;                 assign ID_S_32a32f8d_795a5f17_E[ 14]  =  5'd31;                 assign ID_S_32a32f8d_795a5f17_E[ 15]  =  5'd27;                 assign ID_S_32a32f8d_795a5f17_E[ 16]  =  5'd19;                 assign ID_S_32a32f8d_795a5f17_E[ 17]  =  5'd3;                 assign ID_S_32a32f8d_795a5f17_E[ 18]  =  5'd6;                 assign ID_S_32a32f8d_795a5f17_E[ 19]  =  5'd12;                 assign ID_S_32a32f8d_795a5f17_E[ 20]  =  5'd24;                 assign ID_S_32a32f8d_795a5f17_E[ 21]  =  5'd21;                 assign ID_S_32a32f8d_795a5f17_E[ 22]  =  5'd15;                 assign ID_S_32a32f8d_795a5f17_E[ 23]  =  5'd30;                 assign ID_S_32a32f8d_795a5f17_E[ 24]  =  5'd25;                 assign ID_S_32a32f8d_795a5f17_E[ 25]  =  5'd23;                 assign ID_S_32a32f8d_795a5f17_E[ 26]  =  5'd11;                 assign ID_S_32a32f8d_795a5f17_E[ 27]  =  5'd22;                 assign ID_S_32a32f8d_795a5f17_E[ 28]  =  5'd9;                 assign ID_S_32a32f8d_795a5f17_E[ 29]  =  5'd18;                 assign ID_S_32a32f8d_795a5f17_E[ 30]  =  5'd1;            end         4'd6:            begin                  assign ID_S_32a32f8d_795a5f17_E[  0]  =  6'd2;                 assign ID_S_32a32f8d_795a5f17_E[  1]  =  6'd4;                 assign ID_S_32a32f8d_795a5f17_E[  2]  =  6'd8;                 assign ID_S_32a32f8d_795a5f17_E[  3]  =  6'd16;                  assign ID_S_32a32f8d_795a5f17_E[  4]  =  6'd32;                 assign ID_S_32a32f8d_795a5f17_E[  5]  =  6'd3;                 assign ID_S_32a32f8d_795a5f17_E[  6]  =  6'd6;                 assign ID_S_32a32f8d_795a5f17_E[  7]  =  6'd12;                  assign ID_S_32a32f8d_795a5f17_E[  8]  =  6'd24;                 assign ID_S_32a32f8d_795a5f17_E[  9]  =  6'd48;                 assign ID_S_32a32f8d_795a5f17_E[ 10]  =  6'd35;                 assign ID_S_32a32f8d_795a5f17_E[ 11]  =  6'd5;                  assign ID_S_32a32f8d_795a5f17_E[ 12]  =  6'd10;                 assign ID_S_32a32f8d_795a5f17_E[ 13]  =  6'd20;                 assign ID_S_32a32f8d_795a5f17_E[ 14]  =  6'd40;                 assign ID_S_32a32f8d_795a5f17_E[ 15]  =  6'd19;                   assign ID_S_32a32f8d_795a5f17_E[ 16]  =  6'd38;                 assign ID_S_32a32f8d_795a5f17_E[ 17]  =  6'd15;                 assign ID_S_32a32f8d_795a5f17_E[ 18]  =  6'd30;                 assign ID_S_32a32f8d_795a5f17_E[ 19]  =  6'd60;                 assign ID_S_32a32f8d_795a5f17_E[ 20]  =  6'd59;                 assign ID_S_32a32f8d_795a5f17_E[ 21]  =  6'd53;                 assign ID_S_32a32f8d_795a5f17_E[ 22]  =  6'd41;                 assign ID_S_32a32f8d_795a5f17_E[ 23]  =  6'd17;                 assign ID_S_32a32f8d_795a5f17_E[ 24]  =  6'd34;                 assign ID_S_32a32f8d_795a5f17_E[ 25]  =  6'd7;                 assign ID_S_32a32f8d_795a5f17_E[ 26]  =  6'd14;                 assign ID_S_32a32f8d_795a5f17_E[ 27]  =  6'd28;                 assign ID_S_32a32f8d_795a5f17_E[ 28]  =  6'd56;                 assign ID_S_32a32f8d_795a5f17_E[ 29]  =  6'd51;                 assign ID_S_32a32f8d_795a5f17_E[ 30]  =  6'd37;                 assign ID_S_32a32f8d_795a5f17_E[ 31]  =  6'd9;                  assign ID_S_32a32f8d_795a5f17_E[ 32]  =  6'd18;                 assign ID_S_32a32f8d_795a5f17_E[ 33]  =  6'd36;                 assign ID_S_32a32f8d_795a5f17_E[ 34]  =  6'd11;                 assign ID_S_32a32f8d_795a5f17_E[ 35]  =  6'd22;                 assign ID_S_32a32f8d_795a5f17_E[ 36]  =  6'd44;                 assign ID_S_32a32f8d_795a5f17_E[ 37]  =  6'd27;                 assign ID_S_32a32f8d_795a5f17_E[ 38]  =  6'd54;                 assign ID_S_32a32f8d_795a5f17_E[ 39]  =  6'd47;                 assign ID_S_32a32f8d_795a5f17_E[ 40]  =  6'd29;                 assign ID_S_32a32f8d_795a5f17_E[ 41]  =  6'd58;                 assign ID_S_32a32f8d_795a5f17_E[ 42]  =  6'd55;                 assign ID_S_32a32f8d_795a5f17_E[ 43]  =  6'd45;                 assign ID_S_32a32f8d_795a5f17_E[ 44]  =  6'd25;                 assign ID_S_32a32f8d_795a5f17_E[ 45]  =  6'd50;                 assign ID_S_32a32f8d_795a5f17_E[ 46]  =  6'd39;                 assign ID_S_32a32f8d_795a5f17_E[ 47]  =  6'd13;                 assign ID_S_32a32f8d_795a5f17_E[ 48]  =  6'd26;                 assign ID_S_32a32f8d_795a5f17_E[ 49]  =  6'd52;                 assign ID_S_32a32f8d_795a5f17_E[ 50]  =  6'd43;                 assign ID_S_32a32f8d_795a5f17_E[ 51]  =  6'd21;                 assign ID_S_32a32f8d_795a5f17_E[ 52]  =  6'd42;                 assign ID_S_32a32f8d_795a5f17_E[ 53]  =  6'd23;                 assign ID_S_32a32f8d_795a5f17_E[ 54]  =  6'd46;                 assign ID_S_32a32f8d_795a5f17_E[ 55]  =  6'd31;                 assign ID_S_32a32f8d_795a5f17_E[ 56]  =  6'd62;                 assign ID_S_32a32f8d_795a5f17_E[ 57]  =  6'd63;                 assign ID_S_32a32f8d_795a5f17_E[ 58]  =  6'd61;                 assign ID_S_32a32f8d_795a5f17_E[ 59]  =  6'd57;                 assign ID_S_32a32f8d_795a5f17_E[ 60]  =  6'd49;                 assign ID_S_32a32f8d_795a5f17_E[ 61]  =  6'd33;                 assign ID_S_32a32f8d_795a5f17_E[ 62]  =  6'd1;            end         4'd7:            begin               assign ID_S_32a32f8d_795a5f17_E[  0] = 7'd2;                 assign ID_S_32a32f8d_795a5f17_E[  1] = 7'd4;                assign ID_S_32a32f8d_795a5f17_E[  2] = 7'd8;                assign ID_S_32a32f8d_795a5f17_E[  3] = 7'd16;              assign ID_S_32a32f8d_795a5f17_E[  4] = 7'd32;              assign ID_S_32a32f8d_795a5f17_E[  5] = 7'd64;              assign ID_S_32a32f8d_795a5f17_E[  6] = 7'd9;              assign ID_S_32a32f8d_795a5f17_E[  7] = 7'd18;              assign ID_S_32a32f8d_795a5f17_E[  8] = 7'd36;              assign ID_S_32a32f8d_795a5f17_E[  9] = 7'd72;              assign ID_S_32a32f8d_795a5f17_E[ 10] = 7'd25;              assign ID_S_32a32f8d_795a5f17_E[ 11] = 7'd50;              assign ID_S_32a32f8d_795a5f17_E[ 12] = 7'd100;              assign ID_S_32a32f8d_795a5f17_E[ 13] = 7'd65;              assign ID_S_32a32f8d_795a5f17_E[ 14] = 7'd11;              assign ID_S_32a32f8d_795a5f17_E[ 15] = 7'd22;              assign ID_S_32a32f8d_795a5f17_E[ 16] = 7'd44;              assign ID_S_32a32f8d_795a5f17_E[ 17] = 7'd88;              assign ID_S_32a32f8d_795a5f17_E[ 18] = 7'd57;              assign ID_S_32a32f8d_795a5f17_E[ 19] = 7'd114;              assign ID_S_32a32f8d_795a5f17_E[ 20] = 7'd109;              assign ID_S_32a32f8d_795a5f17_E[ 21] = 7'd83;              assign ID_S_32a32f8d_795a5f17_E[ 22] = 7'd47;              assign ID_S_32a32f8d_795a5f17_E[ 23] = 7'd94;              assign ID_S_32a32f8d_795a5f17_E[ 24] = 7'd53;              assign ID_S_32a32f8d_795a5f17_E[ 25] = 7'd106;              assign ID_S_32a32f8d_795a5f17_E[ 26] = 7'd93;              assign ID_S_32a32f8d_795a5f17_E[ 27] = 7'd51;              assign ID_S_32a32f8d_795a5f17_E[ 28] = 7'd102;              assign ID_S_32a32f8d_795a5f17_E[ 29] = 7'd69;              assign ID_S_32a32f8d_795a5f17_E[ 30] = 7'd3;              assign ID_S_32a32f8d_795a5f17_E[ 31] = 7'd6;              assign ID_S_32a32f8d_795a5f17_E[ 32] = 7'd12;              assign ID_S_32a32f8d_795a5f17_E[ 33] = 7'd24;              assign ID_S_32a32f8d_795a5f17_E[ 34] = 7'd48;              assign ID_S_32a32f8d_795a5f17_E[ 35] = 7'd96;              assign ID_S_32a32f8d_795a5f17_E[ 36] = 7'd73;              assign ID_S_32a32f8d_795a5f17_E[ 37] = 7'd27;              assign ID_S_32a32f8d_795a5f17_E[ 38] = 7'd54;              assign ID_S_32a32f8d_795a5f17_E[ 39] = 7'd108;              assign ID_S_32a32f8d_795a5f17_E[ 40] = 7'd81;              assign ID_S_32a32f8d_795a5f17_E[ 41] = 7'd43;              assign ID_S_32a32f8d_795a5f17_E[ 42] = 7'd86;              assign ID_S_32a32f8d_795a5f17_E[ 43] = 7'd37;              assign ID_S_32a32f8d_795a5f17_E[ 44] = 7'd74;              assign ID_S_32a32f8d_795a5f17_E[ 45] = 7'd29;              assign ID_S_32a32f8d_795a5f17_E[ 46] = 7'd58;              assign ID_S_32a32f8d_795a5f17_E[ 47] = 7'd116;              assign ID_S_32a32f8d_795a5f17_E[ 48] = 7'd97;              assign ID_S_32a32f8d_795a5f17_E[ 49] = 7'd75;              assign ID_S_32a32f8d_795a5f17_E[ 50] = 7'd31;              assign ID_S_32a32f8d_795a5f17_E[ 51] = 7'd62;              assign ID_S_32a32f8d_795a5f17_E[ 52] = 7'd124;              assign ID_S_32a32f8d_795a5f17_E[ 53] = 7'd113;              assign ID_S_32a32f8d_795a5f17_E[ 54] = 7'd107;              assign ID_S_32a32f8d_795a5f17_E[ 55] = 7'd95;              assign ID_S_32a32f8d_795a5f17_E[ 56] = 7'd55;              assign ID_S_32a32f8d_795a5f17_E[ 57] = 7'd110;              assign ID_S_32a32f8d_795a5f17_E[ 58] = 7'd85;              assign ID_S_32a32f8d_795a5f17_E[ 59] = 7'd35;              assign ID_S_32a32f8d_795a5f17_E[ 60] = 7'd70;              assign ID_S_32a32f8d_795a5f17_E[ 61] = 7'd5;              assign ID_S_32a32f8d_795a5f17_E[ 62] = 7'd10;              assign ID_S_32a32f8d_795a5f17_E[ 63] = 7'd20;              assign ID_S_32a32f8d_795a5f17_E[ 64] = 7'd40;              assign ID_S_32a32f8d_795a5f17_E[ 65] = 7'd80;              assign ID_S_32a32f8d_795a5f17_E[ 66] = 7'd41;              assign ID_S_32a32f8d_795a5f17_E[ 67] = 7'd82;              assign ID_S_32a32f8d_795a5f17_E[ 68] = 7'd45;              assign ID_S_32a32f8d_795a5f17_E[ 69] = 7'd90;              assign ID_S_32a32f8d_795a5f17_E[ 70] = 7'd61;              assign ID_S_32a32f8d_795a5f17_E[ 71] = 7'd122;              assign ID_S_32a32f8d_795a5f17_E[ 72] = 7'd125;              assign ID_S_32a32f8d_795a5f17_E[ 73] = 7'd115;              assign ID_S_32a32f8d_795a5f17_E[ 74] = 7'd111;              assign ID_S_32a32f8d_795a5f17_E[ 75] = 7'd87;              assign ID_S_32a32f8d_795a5f17_E[ 76] = 7'd39;              assign ID_S_32a32f8d_795a5f17_E[ 77] = 7'd78;              assign ID_S_32a32f8d_795a5f17_E[ 78] = 7'd21;              assign ID_S_32a32f8d_795a5f17_E[ 79] = 7'd42;              assign ID_S_32a32f8d_795a5f17_E[ 80] = 7'd84;              assign ID_S_32a32f8d_795a5f17_E[ 81] = 7'd33;              assign ID_S_32a32f8d_795a5f17_E[ 82] = 7'd66;              assign ID_S_32a32f8d_795a5f17_E[ 83] = 7'd13;              assign ID_S_32a32f8d_795a5f17_E[ 84] = 7'd26;              assign ID_S_32a32f8d_795a5f17_E[ 85] = 7'd52;              assign ID_S_32a32f8d_795a5f17_E[ 86] = 7'd104;              assign ID_S_32a32f8d_795a5f17_E[ 87] = 7'd89;              assign ID_S_32a32f8d_795a5f17_E[ 88] = 7'd59;              assign ID_S_32a32f8d_795a5f17_E[ 89] = 7'd118;              assign ID_S_32a32f8d_795a5f17_E[ 90] = 7'd101;              assign ID_S_32a32f8d_795a5f17_E[ 91] = 7'd67;              assign ID_S_32a32f8d_795a5f17_E[ 92] = 7'd15;              assign ID_S_32a32f8d_795a5f17_E[ 93] = 7'd30;              assign ID_S_32a32f8d_795a5f17_E[ 94] = 7'd60;              assign ID_S_32a32f8d_795a5f17_E[ 95] = 7'd120;              assign ID_S_32a32f8d_795a5f17_E[ 96] = 7'd121;              assign ID_S_32a32f8d_795a5f17_E[ 97] = 7'd123;              assign ID_S_32a32f8d_795a5f17_E[ 98] = 7'd127;              assign ID_S_32a32f8d_795a5f17_E[ 99] = 7'd119;              assign ID_S_32a32f8d_795a5f17_E[100] = 7'd103;              assign ID_S_32a32f8d_795a5f17_E[101] = 7'd71;              assign ID_S_32a32f8d_795a5f17_E[102] = 7'd7;              assign ID_S_32a32f8d_795a5f17_E[103] = 7'd14;              assign ID_S_32a32f8d_795a5f17_E[104] = 7'd28;              assign ID_S_32a32f8d_795a5f17_E[105] = 7'd56;              assign ID_S_32a32f8d_795a5f17_E[106] = 7'd112;              assign ID_S_32a32f8d_795a5f17_E[107] = 7'd105;              assign ID_S_32a32f8d_795a5f17_E[108] = 7'd91;              assign ID_S_32a32f8d_795a5f17_E[109] = 7'd63;              assign ID_S_32a32f8d_795a5f17_E[110] = 7'd126;              assign ID_S_32a32f8d_795a5f17_E[111] = 7'd117;              assign ID_S_32a32f8d_795a5f17_E[112] = 7'd99;              assign ID_S_32a32f8d_795a5f17_E[113] = 7'd79;              assign ID_S_32a32f8d_795a5f17_E[114] = 7'd23;              assign ID_S_32a32f8d_795a5f17_E[115] = 7'd46;              assign ID_S_32a32f8d_795a5f17_E[116] = 7'd92;              assign ID_S_32a32f8d_795a5f17_E[117] = 7'd49;              assign ID_S_32a32f8d_795a5f17_E[118] = 7'd98;              assign ID_S_32a32f8d_795a5f17_E[119] = 7'd77;              assign ID_S_32a32f8d_795a5f17_E[120] = 7'd19;              assign ID_S_32a32f8d_795a5f17_E[121] = 7'd38;              assign ID_S_32a32f8d_795a5f17_E[122] = 7'd76;              assign ID_S_32a32f8d_795a5f17_E[123] = 7'd17;              assign ID_S_32a32f8d_795a5f17_E[124] = 7'd34;              assign ID_S_32a32f8d_795a5f17_E[125] = 7'd68;              assign ID_S_32a32f8d_795a5f17_E[126] = 7'd1;                                            end         4'd8:             begin                  assign ID_S_32a32f8d_795a5f17_E[  0] = 8'd2;                 assign ID_S_32a32f8d_795a5f17_E[  1] = 8'd4;                                 assign ID_S_32a32f8d_795a5f17_E[  2] = 8'd8;                 assign ID_S_32a32f8d_795a5f17_E[  3] = 8'd16;                 assign ID_S_32a32f8d_795a5f17_E[  4] = 8'd32;                 assign ID_S_32a32f8d_795a5f17_E[  5] = 8'd64;                 assign ID_S_32a32f8d_795a5f17_E[  6] = 8'd128;                 assign ID_S_32a32f8d_795a5f17_E[  7] = 8'd29;                 assign ID_S_32a32f8d_795a5f17_E[  8] = 8'd58;                 assign ID_S_32a32f8d_795a5f17_E[  9] = 8'd116;                 assign ID_S_32a32f8d_795a5f17_E[ 10] = 8'd232;                 assign ID_S_32a32f8d_795a5f17_E[ 11] = 8'd205;                 assign ID_S_32a32f8d_795a5f17_E[ 12] = 8'd135;                 assign ID_S_32a32f8d_795a5f17_E[ 13] = 8'd19;                 assign ID_S_32a32f8d_795a5f17_E[ 14] = 8'd38;                 assign ID_S_32a32f8d_795a5f17_E[ 15] = 8'd76;                 assign ID_S_32a32f8d_795a5f17_E[ 16] = 8'd152;                 assign ID_S_32a32f8d_795a5f17_E[ 17] = 8'd45;                 assign ID_S_32a32f8d_795a5f17_E[ 18] = 8'd90;                 assign ID_S_32a32f8d_795a5f17_E[ 19] = 8'd180;                 assign ID_S_32a32f8d_795a5f17_E[ 20] = 8'd117;                 assign ID_S_32a32f8d_795a5f17_E[ 21] = 8'd234;                 assign ID_S_32a32f8d_795a5f17_E[ 22] = 8'd201;                 assign ID_S_32a32f8d_795a5f17_E[ 23] = 8'd143;                 assign ID_S_32a32f8d_795a5f17_E[ 24] = 8'd3;                 assign ID_S_32a32f8d_795a5f17_E[ 25] = 8'd6;                 assign ID_S_32a32f8d_795a5f17_E[ 26] = 8'd12;                 assign ID_S_32a32f8d_795a5f17_E[ 27] = 8'd24;                 assign ID_S_32a32f8d_795a5f17_E[ 28] = 8'd48;                 assign ID_S_32a32f8d_795a5f17_E[ 29] = 8'd96;                 assign ID_S_32a32f8d_795a5f17_E[ 30] = 8'd192;                 assign ID_S_32a32f8d_795a5f17_E[ 31] = 8'd157;                 assign ID_S_32a32f8d_795a5f17_E[ 32] = 8'd39;                 assign ID_S_32a32f8d_795a5f17_E[ 33] = 8'd78;                 assign ID_S_32a32f8d_795a5f17_E[ 34] = 8'd156;                 assign ID_S_32a32f8d_795a5f17_E[ 35] = 8'd37;                 assign ID_S_32a32f8d_795a5f17_E[ 36] = 8'd74;                 assign ID_S_32a32f8d_795a5f17_E[ 37] = 8'd148;                 assign ID_S_32a32f8d_795a5f17_E[ 38] = 8'd53;                 assign ID_S_32a32f8d_795a5f17_E[ 39] = 8'd106;                 assign ID_S_32a32f8d_795a5f17_E[ 40] = 8'd212;                 assign ID_S_32a32f8d_795a5f17_E[ 41] = 8'd181;                 assign ID_S_32a32f8d_795a5f17_E[ 42] = 8'd119;                 assign ID_S_32a32f8d_795a5f17_E[ 43] = 8'd238;                 assign ID_S_32a32f8d_795a5f17_E[ 44] = 8'd193;                 assign ID_S_32a32f8d_795a5f17_E[ 45] = 8'd159;                 assign ID_S_32a32f8d_795a5f17_E[ 46] = 8'd35;                 assign ID_S_32a32f8d_795a5f17_E[ 47] = 8'd70;                 assign ID_S_32a32f8d_795a5f17_E[ 48] = 8'd140;                 assign ID_S_32a32f8d_795a5f17_E[ 49] = 8'd5;                 assign ID_S_32a32f8d_795a5f17_E[ 50] = 8'd10;                 assign ID_S_32a32f8d_795a5f17_E[ 51] = 8'd20;                 assign ID_S_32a32f8d_795a5f17_E[ 52] = 8'd40;                 assign ID_S_32a32f8d_795a5f17_E[ 53] = 8'd80;                 assign ID_S_32a32f8d_795a5f17_E[ 54] = 8'd160;                 assign ID_S_32a32f8d_795a5f17_E[ 55] = 8'd93;                 assign ID_S_32a32f8d_795a5f17_E[ 56] = 8'd186;                 assign ID_S_32a32f8d_795a5f17_E[ 57] = 8'd105;                 assign ID_S_32a32f8d_795a5f17_E[ 58] = 8'd210;                 assign ID_S_32a32f8d_795a5f17_E[ 59] = 8'd185;                 assign ID_S_32a32f8d_795a5f17_E[ 60] = 8'd111;                 assign ID_S_32a32f8d_795a5f17_E[ 61] = 8'd222;                 assign ID_S_32a32f8d_795a5f17_E[ 62] = 8'd161;                 assign ID_S_32a32f8d_795a5f17_E[ 63] = 8'd95;                 assign ID_S_32a32f8d_795a5f17_E[ 64] = 8'd190;                 assign ID_S_32a32f8d_795a5f17_E[ 65] = 8'd97;                 assign ID_S_32a32f8d_795a5f17_E[ 66] = 8'd194;                 assign ID_S_32a32f8d_795a5f17_E[ 67] = 8'd153;                 assign ID_S_32a32f8d_795a5f17_E[ 68] = 8'd47;                 assign ID_S_32a32f8d_795a5f17_E[ 69] = 8'd94;                 assign ID_S_32a32f8d_795a5f17_E[ 70] = 8'd188;                 assign ID_S_32a32f8d_795a5f17_E[ 71] = 8'd101;                 assign ID_S_32a32f8d_795a5f17_E[ 72] = 8'd202;                 assign ID_S_32a32f8d_795a5f17_E[ 73] = 8'd137;                 assign ID_S_32a32f8d_795a5f17_E[ 74] = 8'd15;                 assign ID_S_32a32f8d_795a5f17_E[ 75] = 8'd30;                 assign ID_S_32a32f8d_795a5f17_E[ 76] = 8'd60;                 assign ID_S_32a32f8d_795a5f17_E[ 77] = 8'd120;                 assign ID_S_32a32f8d_795a5f17_E[ 78] = 8'd240;                 assign ID_S_32a32f8d_795a5f17_E[ 79] = 8'd253;                 assign ID_S_32a32f8d_795a5f17_E[ 80] = 8'd231;                 assign ID_S_32a32f8d_795a5f17_E[ 81] = 8'd211;                 assign ID_S_32a32f8d_795a5f17_E[ 82] = 8'd187;                 assign ID_S_32a32f8d_795a5f17_E[ 83] = 8'd107;                 assign ID_S_32a32f8d_795a5f17_E[ 84] = 8'd214;                 assign ID_S_32a32f8d_795a5f17_E[ 85] = 8'd177;                 assign ID_S_32a32f8d_795a5f17_E[ 86] = 8'd127;                 assign ID_S_32a32f8d_795a5f17_E[ 87] = 8'd254;                 assign ID_S_32a32f8d_795a5f17_E[ 88] = 8'd225;                 assign ID_S_32a32f8d_795a5f17_E[ 89] = 8'd223;                 assign ID_S_32a32f8d_795a5f17_E[ 90] = 8'd163;                 assign ID_S_32a32f8d_795a5f17_E[ 91] = 8'd91;                 assign ID_S_32a32f8d_795a5f17_E[ 92] = 8'd182;                 assign ID_S_32a32f8d_795a5f17_E[ 93] = 8'd113;                 assign ID_S_32a32f8d_795a5f17_E[ 94] = 8'd226;                 assign ID_S_32a32f8d_795a5f17_E[ 95] = 8'd217;                 assign ID_S_32a32f8d_795a5f17_E[ 96] = 8'd175;                 assign ID_S_32a32f8d_795a5f17_E[ 97] = 8'd67;                 assign ID_S_32a32f8d_795a5f17_E[ 98] = 8'd134;                 assign ID_S_32a32f8d_795a5f17_E[ 99] = 8'd17;                 assign ID_S_32a32f8d_795a5f17_E[100] = 8'd34;                 assign ID_S_32a32f8d_795a5f17_E[101] = 8'd68;                 assign ID_S_32a32f8d_795a5f17_E[102] = 8'd136;                 assign ID_S_32a32f8d_795a5f17_E[103] = 8'd13;                 assign ID_S_32a32f8d_795a5f17_E[104] = 8'd26;                 assign ID_S_32a32f8d_795a5f17_E[105] = 8'd52;                 assign ID_S_32a32f8d_795a5f17_E[106] = 8'd104;                 assign ID_S_32a32f8d_795a5f17_E[107] = 8'd208;                 assign ID_S_32a32f8d_795a5f17_E[108] = 8'd189;                 assign ID_S_32a32f8d_795a5f17_E[109] = 8'd103;                 assign ID_S_32a32f8d_795a5f17_E[110] = 8'd206;                 assign ID_S_32a32f8d_795a5f17_E[111] = 8'd129;                 assign ID_S_32a32f8d_795a5f17_E[112] = 8'd31;                 assign ID_S_32a32f8d_795a5f17_E[113] = 8'd62;                 assign ID_S_32a32f8d_795a5f17_E[114] = 8'd124;                 assign ID_S_32a32f8d_795a5f17_E[115] = 8'd248;                 assign ID_S_32a32f8d_795a5f17_E[116] = 8'd237;                 assign ID_S_32a32f8d_795a5f17_E[117] = 8'd199;                 assign ID_S_32a32f8d_795a5f17_E[118] = 8'd147;                 assign ID_S_32a32f8d_795a5f17_E[119] = 8'd59;                 assign ID_S_32a32f8d_795a5f17_E[120] = 8'd118;                 assign ID_S_32a32f8d_795a5f17_E[121] = 8'd236;                 assign ID_S_32a32f8d_795a5f17_E[122] = 8'd197;                 assign ID_S_32a32f8d_795a5f17_E[123] = 8'd151;                 assign ID_S_32a32f8d_795a5f17_E[124] = 8'd51;                 assign ID_S_32a32f8d_795a5f17_E[125] = 8'd102;                 assign ID_S_32a32f8d_795a5f17_E[126] = 8'd204;                 assign ID_S_32a32f8d_795a5f17_E[127] = 8'd133;                 assign ID_S_32a32f8d_795a5f17_E[128] = 8'd23;                 assign ID_S_32a32f8d_795a5f17_E[129] = 8'd46;                 assign ID_S_32a32f8d_795a5f17_E[130] = 8'd92;                 assign ID_S_32a32f8d_795a5f17_E[131] = 8'd184;                 assign ID_S_32a32f8d_795a5f17_E[132] = 8'd109;                 assign ID_S_32a32f8d_795a5f17_E[133] = 8'd218;                                 assign ID_S_32a32f8d_795a5f17_E[134] = 8'd169;                                 assign ID_S_32a32f8d_795a5f17_E[135] = 8'd79;                                 assign ID_S_32a32f8d_795a5f17_E[136] = 8'd158;                                 assign ID_S_32a32f8d_795a5f17_E[137] = 8'd33;                                 assign ID_S_32a32f8d_795a5f17_E[138] = 8'd66;                                 assign ID_S_32a32f8d_795a5f17_E[139] = 8'd132;                                 assign ID_S_32a32f8d_795a5f17_E[140] = 8'd21;                                 assign ID_S_32a32f8d_795a5f17_E[141] = 8'd42;                                 assign ID_S_32a32f8d_795a5f17_E[142] = 8'd84;                                 assign ID_S_32a32f8d_795a5f17_E[143] = 8'd168;                                 assign ID_S_32a32f8d_795a5f17_E[144] = 8'd77;                                 assign ID_S_32a32f8d_795a5f17_E[145] = 8'd154;                                 assign ID_S_32a32f8d_795a5f17_E[146] = 8'd41;                                 assign ID_S_32a32f8d_795a5f17_E[147] = 8'd82;                                 assign ID_S_32a32f8d_795a5f17_E[148] = 8'd164;                                 assign ID_S_32a32f8d_795a5f17_E[149] = 8'd85;                                 assign ID_S_32a32f8d_795a5f17_E[150] = 8'd170;                                 assign ID_S_32a32f8d_795a5f17_E[151] = 8'd73;                                 assign ID_S_32a32f8d_795a5f17_E[152] = 8'd146;                                 assign ID_S_32a32f8d_795a5f17_E[153] = 8'd57;                                 assign ID_S_32a32f8d_795a5f17_E[154] = 8'd114;                                 assign ID_S_32a32f8d_795a5f17_E[155] = 8'd228;                                 assign ID_S_32a32f8d_795a5f17_E[156] = 8'd213;                                 assign ID_S_32a32f8d_795a5f17_E[157] = 8'd183;                                 assign ID_S_32a32f8d_795a5f17_E[158] = 8'd115;                                 assign ID_S_32a32f8d_795a5f17_E[159] = 8'd230;                                 assign ID_S_32a32f8d_795a5f17_E[160] = 8'd209;                                 assign ID_S_32a32f8d_795a5f17_E[161] = 8'd191;                                 assign ID_S_32a32f8d_795a5f17_E[162] = 8'd99;                                 assign ID_S_32a32f8d_795a5f17_E[163] = 8'd198;                                 assign ID_S_32a32f8d_795a5f17_E[164] = 8'd145;                                 assign ID_S_32a32f8d_795a5f17_E[165] = 8'd63;                                 assign ID_S_32a32f8d_795a5f17_E[166] = 8'd126;                 assign ID_S_32a32f8d_795a5f17_E[167] = 8'd252;                 assign ID_S_32a32f8d_795a5f17_E[168] = 8'd229;                 assign ID_S_32a32f8d_795a5f17_E[169] = 8'd215;                 assign ID_S_32a32f8d_795a5f17_E[170] = 8'd179;                 assign ID_S_32a32f8d_795a5f17_E[171] = 8'd123;                 assign ID_S_32a32f8d_795a5f17_E[172] = 8'd246;                 assign ID_S_32a32f8d_795a5f17_E[173] = 8'd241;                 assign ID_S_32a32f8d_795a5f17_E[174] = 8'd255;                 assign ID_S_32a32f8d_795a5f17_E[175] = 8'd227;                 assign ID_S_32a32f8d_795a5f17_E[176] = 8'd219;                 assign ID_S_32a32f8d_795a5f17_E[177] = 8'd171;                 assign ID_S_32a32f8d_795a5f17_E[178] = 8'd75;                 assign ID_S_32a32f8d_795a5f17_E[179] = 8'd150;                 assign ID_S_32a32f8d_795a5f17_E[180] = 8'd49;                 assign ID_S_32a32f8d_795a5f17_E[181] = 8'd98;                 assign ID_S_32a32f8d_795a5f17_E[182] = 8'd196;                 assign ID_S_32a32f8d_795a5f17_E[183] = 8'd149;                 assign ID_S_32a32f8d_795a5f17_E[184] = 8'd55;                 assign ID_S_32a32f8d_795a5f17_E[185] = 8'd110;                 assign ID_S_32a32f8d_795a5f17_E[186] = 8'd220;                 assign ID_S_32a32f8d_795a5f17_E[187] = 8'd165;                 assign ID_S_32a32f8d_795a5f17_E[188] = 8'd87;                 assign ID_S_32a32f8d_795a5f17_E[189] = 8'd174;                 assign ID_S_32a32f8d_795a5f17_E[190] = 8'd65;                 assign ID_S_32a32f8d_795a5f17_E[191] = 8'd130;                 assign ID_S_32a32f8d_795a5f17_E[192] = 8'd25;                 assign ID_S_32a32f8d_795a5f17_E[193] = 8'd50;                 assign ID_S_32a32f8d_795a5f17_E[194] = 8'd100;                 assign ID_S_32a32f8d_795a5f17_E[195] = 8'd200;                 assign ID_S_32a32f8d_795a5f17_E[196] = 8'd141;                 assign ID_S_32a32f8d_795a5f17_E[197] = 8'd7;                 assign ID_S_32a32f8d_795a5f17_E[198] = 8'd14;                 assign ID_S_32a32f8d_795a5f17_E[199] = 8'd28;                 assign ID_S_32a32f8d_795a5f17_E[200] = 8'd56;                 assign ID_S_32a32f8d_795a5f17_E[201] = 8'd112;                 assign ID_S_32a32f8d_795a5f17_E[202] = 8'd224;                 assign ID_S_32a32f8d_795a5f17_E[203] = 8'd221;                 assign ID_S_32a32f8d_795a5f17_E[204] = 8'd167;                 assign ID_S_32a32f8d_795a5f17_E[205] = 8'd83;                 assign ID_S_32a32f8d_795a5f17_E[206] = 8'd166;                 assign ID_S_32a32f8d_795a5f17_E[207] = 8'd81;                 assign ID_S_32a32f8d_795a5f17_E[208] = 8'd62;                 assign ID_S_32a32f8d_795a5f17_E[209] = 8'd89;                 assign ID_S_32a32f8d_795a5f17_E[210] = 8'd178;                 assign ID_S_32a32f8d_795a5f17_E[211] = 8'd121;                 assign ID_S_32a32f8d_795a5f17_E[212] = 8'd242;                 assign ID_S_32a32f8d_795a5f17_E[213] = 8'd249;                 assign ID_S_32a32f8d_795a5f17_E[214] = 8'd239;                 assign ID_S_32a32f8d_795a5f17_E[215] = 8'd195;                 assign ID_S_32a32f8d_795a5f17_E[216] = 8'd155;                 assign ID_S_32a32f8d_795a5f17_E[217] = 8'd43;                 assign ID_S_32a32f8d_795a5f17_E[218] = 8'd86;                 assign ID_S_32a32f8d_795a5f17_E[219] = 8'd172;                 assign ID_S_32a32f8d_795a5f17_E[220] = 8'd69;                 assign ID_S_32a32f8d_795a5f17_E[221] = 8'd138;                 assign ID_S_32a32f8d_795a5f17_E[222] = 8'd9;                 assign ID_S_32a32f8d_795a5f17_E[223] = 8'd18;                 assign ID_S_32a32f8d_795a5f17_E[224] = 8'd36;                 assign ID_S_32a32f8d_795a5f17_E[225] = 8'd72;                 assign ID_S_32a32f8d_795a5f17_E[226] = 8'd144;                 assign ID_S_32a32f8d_795a5f17_E[227] = 8'd61;                 assign ID_S_32a32f8d_795a5f17_E[228] = 8'd122;                 assign ID_S_32a32f8d_795a5f17_E[229] = 8'd244;                 assign ID_S_32a32f8d_795a5f17_E[230] = 8'd245;                 assign ID_S_32a32f8d_795a5f17_E[231] = 8'd247;                 assign ID_S_32a32f8d_795a5f17_E[232] = 8'd243;                 assign ID_S_32a32f8d_795a5f17_E[233] = 8'd251;                 assign ID_S_32a32f8d_795a5f17_E[234] = 8'd235;                 assign ID_S_32a32f8d_795a5f17_E[235] = 8'd203;                 assign ID_S_32a32f8d_795a5f17_E[236] = 8'd139;                 assign ID_S_32a32f8d_795a5f17_E[237] = 8'd11;                 assign ID_S_32a32f8d_795a5f17_E[238] = 8'd22;                 assign ID_S_32a32f8d_795a5f17_E[239] = 8'd44;                 assign ID_S_32a32f8d_795a5f17_E[240] = 8'd88;                 assign ID_S_32a32f8d_795a5f17_E[241] = 8'd176;                 assign ID_S_32a32f8d_795a5f17_E[242] = 8'd125;                 assign ID_S_32a32f8d_795a5f17_E[243] = 8'd250;                 assign ID_S_32a32f8d_795a5f17_E[244] = 8'd233;                 assign ID_S_32a32f8d_795a5f17_E[245] = 8'd207;                 assign ID_S_32a32f8d_795a5f17_E[246] = 8'd131;                 assign ID_S_32a32f8d_795a5f17_E[247] = 8'd27;                 assign ID_S_32a32f8d_795a5f17_E[248] = 8'd54;                 assign ID_S_32a32f8d_795a5f17_E[249] = 8'd108;                 assign ID_S_32a32f8d_795a5f17_E[250] = 8'd216;                 assign ID_S_32a32f8d_795a5f17_E[251] = 8'd173;                 assign ID_S_32a32f8d_795a5f17_E[252] = 8'd71;                 assign ID_S_32a32f8d_795a5f17_E[253] = 8'd142;                 assign ID_S_32a32f8d_795a5f17_E[254] = 8'd1  ;                 end                       endcase endgenerate  reg [SYM_BW-1:0]  ID_S_f176c2b_400d4b5a_E[T_NUM-1:0];  wire [SYM_BW-1:0] ID_S_1439373b_2f1ff4ba_E[T_NUM-1:0];  wire [SYM_BW-1:0] ID_S_7c9e683d_1f35ac67_E[T_NUM-1:0];  wire [SYM_BW-1:0] ID_S_71534e04_678b7aad_E;   reg [SYM_BW-1:0] ID_S_526ef0a1_367942f8_E[T_NUM:0];      genvar ID_S_526eca48_36158cfe_E; generate     for(ID_S_526eca48_36158cfe_E = 0;ID_S_526eca48_36158cfe_E <= T_NUM ;ID_S_526eca48_36158cfe_E = ID_S_526eca48_36158cfe_E + 1)     begin         always @(posedge clk or negedge rst_n)         if (!rst_n) begin                         ID_S_526ef0a1_367942f8_E[ID_S_526eca48_36158cfe_E]    <= 8'd0;                     end else if (start) begin                         ID_S_526ef0a1_367942f8_E[ID_S_526eca48_36158cfe_E]    <= lamda[(ID_S_526eca48_36158cfe_E+1) *SYM_BW - 1:ID_S_526eca48_36158cfe_E *SYM_BW]   ;                          end else ;     end endgenerate   genvar ID_S_682d6daf_65285649_E; generate     for(ID_S_682d6daf_65285649_E = 0;ID_S_682d6daf_65285649_E < T_NUM  ;ID_S_682d6daf_65285649_E = ID_S_682d6daf_65285649_E + 1)     begin         case({SYM_BW})             {4'd3}:             begin:gf8mul_dec                 gf8mul_dec   ID_S_636bb82b_1ce12ccd_E( ID_S_f176c2b_400d4b5a_E[ID_S_682d6daf_65285649_E] ,  ID_S_32a32f8d_795a5f17_E[ID_S_682d6daf_65285649_E]     ,  ID_S_1439373b_2f1ff4ba_E[ID_S_682d6daf_65285649_E] );                 gf8mul_dec   ID_S_637dd0ac_1c136950_E( ID_S_f176c2b_400d4b5a_E[ID_S_682d6daf_65285649_E] ,  ID_S_526ef0a1_367942f8_E[ID_S_682d6daf_65285649_E+1] ,  ID_S_7c9e683d_1f35ac67_E[ID_S_682d6daf_65285649_E]   );                     end                                                                                                      {4'd4}:                                                                                                  begin:gf16mul_dec                                                                                            gf16mul_dec  ID_S_636bb82b_1ce12ccd_E( ID_S_f176c2b_400d4b5a_E[ID_S_682d6daf_65285649_E] ,  ID_S_32a32f8d_795a5f17_E[ID_S_682d6daf_65285649_E]     ,  ID_S_1439373b_2f1ff4ba_E[ID_S_682d6daf_65285649_E] );                 gf16mul_dec  ID_S_637dd0ac_1c136950_E( ID_S_f176c2b_400d4b5a_E[ID_S_682d6daf_65285649_E] ,  ID_S_526ef0a1_367942f8_E[ID_S_682d6daf_65285649_E+1] ,  ID_S_7c9e683d_1f35ac67_E[ID_S_682d6daf_65285649_E]   );                     end                                                                                                      {4'd5}:                                                                                                  begin:gf32mul_dec                                                                                            gf32mul_dec  ID_S_636bb82b_1ce12ccd_E( ID_S_f176c2b_400d4b5a_E[ID_S_682d6daf_65285649_E] ,  ID_S_32a32f8d_795a5f17_E[ID_S_682d6daf_65285649_E]     ,  ID_S_1439373b_2f1ff4ba_E[ID_S_682d6daf_65285649_E] );                 gf32mul_dec  ID_S_637dd0ac_1c136950_E( ID_S_f176c2b_400d4b5a_E[ID_S_682d6daf_65285649_E] ,  ID_S_526ef0a1_367942f8_E[ID_S_682d6daf_65285649_E+1] ,  ID_S_7c9e683d_1f35ac67_E[ID_S_682d6daf_65285649_E]   );                     end                                                                                                      {4'd6}:                                                                                                  begin:gf64mul_dec                                                                                            gf64mul_dec  ID_S_636bb82b_1ce12ccd_E( ID_S_f176c2b_400d4b5a_E[ID_S_682d6daf_65285649_E] ,  ID_S_32a32f8d_795a5f17_E[ID_S_682d6daf_65285649_E]     ,  ID_S_1439373b_2f1ff4ba_E[ID_S_682d6daf_65285649_E] );                 gf64mul_dec  ID_S_637dd0ac_1c136950_E( ID_S_f176c2b_400d4b5a_E[ID_S_682d6daf_65285649_E] ,  ID_S_526ef0a1_367942f8_E[ID_S_682d6daf_65285649_E+1] ,  ID_S_7c9e683d_1f35ac67_E[ID_S_682d6daf_65285649_E]   );                     end                                                                                                      {4'd7}:                                                                                                  begin:gf128mul_dec                                                                                           gf128mul_dec ID_S_636bb82b_1ce12ccd_E( ID_S_f176c2b_400d4b5a_E[ID_S_682d6daf_65285649_E] ,  ID_S_32a32f8d_795a5f17_E[ID_S_682d6daf_65285649_E]     ,  ID_S_1439373b_2f1ff4ba_E[ID_S_682d6daf_65285649_E] );                 gf128mul_dec ID_S_637dd0ac_1c136950_E( ID_S_f176c2b_400d4b5a_E[ID_S_682d6daf_65285649_E] ,  ID_S_526ef0a1_367942f8_E[ID_S_682d6daf_65285649_E+1] ,  ID_S_7c9e683d_1f35ac67_E[ID_S_682d6daf_65285649_E]   );                     end                                                                                                                                                                                                               {4'd8}:                                                                                                  begin:gf256mul_dec                                                                                           gf256mul_dec ID_S_636bb82b_1ce12ccd_E( ID_S_f176c2b_400d4b5a_E[ID_S_682d6daf_65285649_E] ,  ID_S_32a32f8d_795a5f17_E[ID_S_682d6daf_65285649_E]     ,  ID_S_1439373b_2f1ff4ba_E[ID_S_682d6daf_65285649_E] );                 gf256mul_dec ID_S_637dd0ac_1c136950_E( ID_S_f176c2b_400d4b5a_E[ID_S_682d6daf_65285649_E] ,  ID_S_526ef0a1_367942f8_E[ID_S_682d6daf_65285649_E+1] ,  ID_S_7c9e683d_1f35ac67_E[ID_S_682d6daf_65285649_E]   );             end         endcase     end endgenerate   generate     case({T_NUM})          
`R_BW'd16:

           begin: ID_S_66c8bbfe_22596c85_E                 assign ID_S_71534e04_678b7aad_E = ID_S_526ef0a1_367942f8_E[0] ^ ID_S_7c9e683d_1f35ac67_E[0] ^ ID_S_7c9e683d_1f35ac67_E[1] ^ ID_S_7c9e683d_1f35ac67_E[2] ^ ID_S_7c9e683d_1f35ac67_E[3] ^ ID_S_7c9e683d_1f35ac67_E[4] ^ ID_S_7c9e683d_1f35ac67_E[5] ^ ID_S_7c9e683d_1f35ac67_E[6] ^ ID_S_7c9e683d_1f35ac67_E[7] ^ ID_S_7c9e683d_1f35ac67_E[8] ^ ID_S_7c9e683d_1f35ac67_E[9] ^ ID_S_7c9e683d_1f35ac67_E[10] ^ ID_S_7c9e683d_1f35ac67_E[11] ^ ID_S_7c9e683d_1f35ac67_E[12] ^ ID_S_7c9e683d_1f35ac67_E[13] ^ ID_S_7c9e683d_1f35ac67_E[14] ^ ID_S_7c9e683d_1f35ac67_E[15];            end         
`R_BW'd8:

           begin : ID_S_7f3c62cf_4f4213db_E                 assign ID_S_71534e04_678b7aad_E = ID_S_526ef0a1_367942f8_E[0] ^ ID_S_7c9e683d_1f35ac67_E[0] ^ ID_S_7c9e683d_1f35ac67_E[1] ^ ID_S_7c9e683d_1f35ac67_E[2] ^ ID_S_7c9e683d_1f35ac67_E[3] ^ ID_S_7c9e683d_1f35ac67_E[4] ^ ID_S_7c9e683d_1f35ac67_E[5] ^ ID_S_7c9e683d_1f35ac67_E[6] ^ ID_S_7c9e683d_1f35ac67_E[7];            end         
`R_BW'd4:

            begin : ID_S_7f3c62cb_4f4213d7_E                 assign ID_S_71534e04_678b7aad_E = ID_S_526ef0a1_367942f8_E[0] ^ ID_S_7c9e683d_1f35ac67_E[0] ^ ID_S_7c9e683d_1f35ac67_E[1] ^ ID_S_7c9e683d_1f35ac67_E[2] ^ ID_S_7c9e683d_1f35ac67_E[3] ;             end         
`R_BW'd2:

            begin : ID_S_7f3c62c9_4f4213d1_E                 assign ID_S_71534e04_678b7aad_E = ID_S_526ef0a1_367942f8_E[0] ^ ID_S_7c9e683d_1f35ac67_E[0] ^ ID_S_7c9e683d_1f35ac67_E[1]  ;             end          
`R_BW'd1:

            begin : ID_S_7f3c62c8_4f4213d2_E                 assign ID_S_71534e04_678b7aad_E = ID_S_526ef0a1_367942f8_E[0] ^ ID_S_7c9e683d_1f35ac67_E[0]  ;             end                 endcase endgenerate       generate     for(ID_S_682d6daf_65285649_E = 0;ID_S_682d6daf_65285649_E < T_NUM  ;ID_S_682d6daf_65285649_E = ID_S_682d6daf_65285649_E + 1)     begin         always @(posedge clk or negedge rst_n)         if (!rst_n)             begin               ID_S_f176c2b_400d4b5a_E[ID_S_682d6daf_65285649_E] <= 0;             end         else if (start)             begin                ID_S_f176c2b_400d4b5a_E[ID_S_682d6daf_65285649_E] <= ID_S_32a32f8d_795a5f17_E[(ID_S_682d6daf_65285649_E+ (ID_S_682d6daf_65285649_E+1)*(ID_S_53b735b7_11413ceb_E)) % (2**SYM_BW - 1)];               end         else if (ID_S_787e79a3_1d07dd47_E)             begin               ID_S_f176c2b_400d4b5a_E[ID_S_682d6daf_65285649_E] <= ID_S_1439373b_2f1ff4ba_E[ID_S_682d6daf_65285649_E];             end         else             ;     end endgenerate    generate     for(ID_S_682d6daf_65285649_E = 0;ID_S_682d6daf_65285649_E < T_NUM  ;ID_S_682d6daf_65285649_E = ID_S_682d6daf_65285649_E + 1)     begin         always @(posedge clk or negedge rst_n)         if (!rst_n)             begin               err_loc[(ID_S_682d6daf_65285649_E+1) *SYM_BW - 1:ID_S_682d6daf_65285649_E *SYM_BW]  <= 0;             end         else if (start)             begin               err_loc[(ID_S_682d6daf_65285649_E+1) *SYM_BW - 1:ID_S_682d6daf_65285649_E *SYM_BW]  <= 0;             end         else if ((ID_S_71534e04_678b7aad_E == 0) && ID_S_787e79a3_1d07dd47_E)             begin                 case(ID_S_6f264d33_7f0e6051_E)                     ID_S_682d6daf_65285649_E: begin err_loc[(ID_S_682d6daf_65285649_E+1) *SYM_BW - 1:ID_S_682d6daf_65285649_E *SYM_BW]  <= ID_S_651d5efd_799ab730_E;   end                 endcase             end         else              ;     end endgenerate   always @(posedge clk or negedge rst_n) if (!rst_n)   ID_S_6f264d33_7f0e6051_E <= 0; else if (start)   ID_S_6f264d33_7f0e6051_E <= 0; else if ((ID_S_71534e04_678b7aad_E == 0) && ID_S_787e79a3_1d07dd47_E)   ID_S_6f264d33_7f0e6051_E <= ID_S_6f264d33_7f0e6051_E + 1;  always @(posedge clk or negedge rst_n) if (!rst_n)     ID_S_651d5efd_799ab730_E <= 0; else if (start)     ID_S_651d5efd_799ab730_E <= 1; else if (ID_S_787e79a3_1d07dd47_E)     ID_S_651d5efd_799ab730_E <= ID_S_651d5efd_799ab730_E + 1; else     ID_S_651d5efd_799ab730_E <= 0;  always @(posedge clk or negedge rst_n) if (!rst_n)     ID_S_787e79a3_1d07dd47_E <= 0; else if (start)      ID_S_787e79a3_1d07dd47_E <= 1;  else if ( ID_S_651d5efd_799ab730_E == N_NUM)     ID_S_787e79a3_1d07dd47_E <= 0; else     ;  always @(posedge clk or negedge rst_n) if (!rst_n)   done <= 0; else if (start )   done <= 0;  else if (ID_S_787e79a3_1d07dd47_E &&  (ID_S_651d5efd_799ab730_E == N_NUM))   done <= 1; else   done <= 0;      endmodule