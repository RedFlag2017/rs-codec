
`timescale 1ns/100ps

module err_value #( parameter [
`SYM_BW_BW -1 :0] SYM_BW = 8,

parameter [8-1:0]  N_NUM = 255, parameter [
`R_BW - 1 :0]  R_NUM = 16,

parameter [
`R_BW - 1 :0]  T_NUM = R_NUM/2

)  (        input clk,        input rst_n,        input start,          input [SYM_BW*(T_NUM+1) - 1:0] lamda,                   input [SYM_BW*(T_NUM) - 1:0] omega,          input [SYM_BW*(T_NUM) - 1:0] err_loc,                        output reg [SYM_BW*(T_NUM) - 1:0] err_val,           output reg [SYM_BW*(T_NUM) - 1:0] err_loc_out,                output reg done        );            localparam ID_S_b8824c0_7ead0f40_E = T_NUM/2;    reg [SYM_BW-1:0] ID_S_678291e7_5121332d_E[T_NUM:0]   ;                 reg [SYM_BW-1:0] ID_S_69e010d1_7dab0633_E[T_NUM - 1:0]   ;  reg [SYM_BW-1:0] ID_S_496ff42e_ba097b9_E[T_NUM - 1:0]   ;     genvar ID_S_526eca48_36158cfe_E; generate     for(ID_S_526eca48_36158cfe_E = 0;ID_S_526eca48_36158cfe_E <= T_NUM ;ID_S_526eca48_36158cfe_E = ID_S_526eca48_36158cfe_E + 1)     begin         always @(posedge clk or negedge rst_n)         if (!rst_n) begin                         ID_S_678291e7_5121332d_E[ID_S_526eca48_36158cfe_E]    <= 8'd0;                     end else if (start) begin             ID_S_678291e7_5121332d_E[ID_S_526eca48_36158cfe_E]    <= lamda[(ID_S_526eca48_36158cfe_E+1) *SYM_BW - 1:ID_S_526eca48_36158cfe_E *SYM_BW]    ;         end else ;     end endgenerate  genvar ID_S_6227abb2_151191de_E; generate     for(ID_S_6227abb2_151191de_E = 0;ID_S_6227abb2_151191de_E < T_NUM   ;ID_S_6227abb2_151191de_E = ID_S_6227abb2_151191de_E + 1)     begin         always @(posedge clk or negedge rst_n)         if (!rst_n) begin                         ID_S_69e010d1_7dab0633_E[ID_S_6227abb2_151191de_E]    <= 8'd0;             ID_S_496ff42e_ba097b9_E[ID_S_6227abb2_151191de_E]    <= 8'd0;         end else if (start) begin             ID_S_69e010d1_7dab0633_E[ID_S_6227abb2_151191de_E]    <= omega[(ID_S_6227abb2_151191de_E+1) *SYM_BW - 1:ID_S_6227abb2_151191de_E *SYM_BW]    ;             ID_S_496ff42e_ba097b9_E[ID_S_6227abb2_151191de_E]    <= err_loc[(ID_S_6227abb2_151191de_E+1) *SYM_BW - 1:ID_S_6227abb2_151191de_E *SYM_BW];         end else ;     end endgenerate     reg [SYM_BW-1:0] ID_S_1cc09e76_634c0c8c_E [T_NUM    :0];       reg [SYM_BW-1:0] ID_S_34d46d67_7fcdf326_E[T_NUM-1  :0];  wire [SYM_BW-1:0] ID_S_1439373b_2f1ff4ba_E[T_NUM:0]; wire [SYM_BW-1:0] ID_S_763fe6b_156a0a07_E[T_NUM-1:0]; reg [8:0] ID_S_651d5efd_799ab730_E;   always @(posedge clk or negedge rst_n) if (!rst_n)   ID_S_651d5efd_799ab730_E <= 0; else if (start)   ID_S_651d5efd_799ab730_E <= 1; else if ((ID_S_651d5efd_799ab730_E < N_NUM ) && ID_S_651d5efd_799ab730_E)   ID_S_651d5efd_799ab730_E <= ID_S_651d5efd_799ab730_E + 1; else    ID_S_651d5efd_799ab730_E <= 0;   wire [SYM_BW-1:0] ID_S_4f622098_66cde942_E [3*16 -1   :0];           generate     case({SYM_BW})          4'd3:            begin                  assign ID_S_4f622098_66cde942_E[0 ]  =  3'd1;                 assign ID_S_4f622098_66cde942_E[1 ]  =  3'd5;                 assign ID_S_4f622098_66cde942_E[2 ]  =  3'd7;                 assign ID_S_4f622098_66cde942_E[3 ]  =  3'd6;                     assign ID_S_4f622098_66cde942_E[4 ]  =  3'd3;                 assign ID_S_4f622098_66cde942_E[5 ]  =  3'd4;            end         4'd4:            begin                  assign ID_S_4f622098_66cde942_E[0 ]  =  4'd1;                 assign ID_S_4f622098_66cde942_E[1 ]  =  4'd9;                 assign ID_S_4f622098_66cde942_E[2 ]  =  4'd13;                 assign ID_S_4f622098_66cde942_E[3 ]  =  4'd15;                                                           assign ID_S_4f622098_66cde942_E[4 ]  =  4'd14;                 assign ID_S_4f622098_66cde942_E[5 ]  =  4'd7;                 assign ID_S_4f622098_66cde942_E[6 ]  =  4'd10;                 assign ID_S_4f622098_66cde942_E[7 ]  =  4'd5;                                                           assign ID_S_4f622098_66cde942_E[8 ]  =  4'd11;                 assign ID_S_4f622098_66cde942_E[9 ]  =  4'd12;                 assign ID_S_4f622098_66cde942_E[10]  =  4'd6;                 assign ID_S_4f622098_66cde942_E[11]  =  4'd3;                            end           4'd5:             begin                  assign ID_S_4f622098_66cde942_E[0 ]  =  5'd1;                 assign ID_S_4f622098_66cde942_E[1 ]  =  5'd18;                 assign ID_S_4f622098_66cde942_E[2 ]  =  5'd9;                 assign ID_S_4f622098_66cde942_E[3 ]  =  5'd22;                  assign ID_S_4f622098_66cde942_E[4 ]  =  5'd11;                 assign ID_S_4f622098_66cde942_E[5 ]  =  5'd23;                 assign ID_S_4f622098_66cde942_E[6 ]  =  5'd25;                 assign ID_S_4f622098_66cde942_E[7 ]  =  5'd30;                  assign ID_S_4f622098_66cde942_E[8 ]  =  5'd15;                 assign ID_S_4f622098_66cde942_E[9 ]  =  5'd21;                 assign ID_S_4f622098_66cde942_E[10]  =  5'd24;                 assign ID_S_4f622098_66cde942_E[11]  =  5'd12;                  assign ID_S_4f622098_66cde942_E[12]  =  5'd6;                 assign ID_S_4f622098_66cde942_E[13]  =  5'd3;                 assign ID_S_4f622098_66cde942_E[14]  =  5'd19;                 assign ID_S_4f622098_66cde942_E[15]  =  5'd27;                                                          assign ID_S_4f622098_66cde942_E[16]  =  5'd31;                                 assign ID_S_4f622098_66cde942_E[17]  =  5'd29;                 assign ID_S_4f622098_66cde942_E[18]  =  5'd28;                 assign ID_S_4f622098_66cde942_E[19]  =  5'd14;                 assign ID_S_4f622098_66cde942_E[20]  =  5'd7;                 assign ID_S_4f622098_66cde942_E[21]  =  5'd17;                 assign ID_S_4f622098_66cde942_E[22]  =  5'd26;                 assign ID_S_4f622098_66cde942_E[23]  =  5'd13;             end              4'd6:             begin                  assign ID_S_4f622098_66cde942_E[0 ]  =  6'd1;                 assign ID_S_4f622098_66cde942_E[1 ]  =  6'd33;                 assign ID_S_4f622098_66cde942_E[2 ]  =  6'd49;                 assign ID_S_4f622098_66cde942_E[3 ]  =  6'd57;                  assign ID_S_4f622098_66cde942_E[4 ]  =  6'd61;                 assign ID_S_4f622098_66cde942_E[5 ]  =  6'd63;                 assign ID_S_4f622098_66cde942_E[6 ]  =  6'd62;                 assign ID_S_4f622098_66cde942_E[7 ]  =  6'd31;                  assign ID_S_4f622098_66cde942_E[8 ]  =  6'd46;                 assign ID_S_4f622098_66cde942_E[9 ]  =  6'd23;                 assign ID_S_4f622098_66cde942_E[10]  =  6'd42;                 assign ID_S_4f622098_66cde942_E[11]  =  6'd21;                  assign ID_S_4f622098_66cde942_E[12]  =  6'd43;                 assign ID_S_4f622098_66cde942_E[13]  =  6'd52;                 assign ID_S_4f622098_66cde942_E[14]  =  6'd26;                 assign ID_S_4f622098_66cde942_E[15]  =  6'd13;                                                          assign ID_S_4f622098_66cde942_E[16]  =  6'd39;                                 assign ID_S_4f622098_66cde942_E[17]  =  6'd50;                 assign ID_S_4f622098_66cde942_E[18]  =  6'd25;                 assign ID_S_4f622098_66cde942_E[19]  =  6'd45;                 assign ID_S_4f622098_66cde942_E[20]  =  6'd55;                 assign ID_S_4f622098_66cde942_E[21]  =  6'd58;                 assign ID_S_4f622098_66cde942_E[22]  =  6'd29;                 assign ID_S_4f622098_66cde942_E[23]  =  6'd47;                 assign ID_S_4f622098_66cde942_E[24]  =  6'd54;                 assign ID_S_4f622098_66cde942_E[25]  =  6'd27;                 assign ID_S_4f622098_66cde942_E[26]  =  6'd44;                 assign ID_S_4f622098_66cde942_E[27]  =  6'd22;                 assign ID_S_4f622098_66cde942_E[28]  =  6'd11;                 assign ID_S_4f622098_66cde942_E[29]  =  6'd36;                 assign ID_S_4f622098_66cde942_E[30]  =  6'd18;                 assign ID_S_4f622098_66cde942_E[31]  =  6'd9;                                                          assign ID_S_4f622098_66cde942_E[32]  =  6'd37;                 assign ID_S_4f622098_66cde942_E[33]  =  6'd51;                 assign ID_S_4f622098_66cde942_E[34]  =  6'd56;                 assign ID_S_4f622098_66cde942_E[35]  =  6'd28;                 assign ID_S_4f622098_66cde942_E[36]  =  6'd14;                 assign ID_S_4f622098_66cde942_E[37]  =  6'd7;                 assign ID_S_4f622098_66cde942_E[38]  =  6'd34;                 assign ID_S_4f622098_66cde942_E[39]  =  6'd17;                 assign ID_S_4f622098_66cde942_E[40]  =  6'd41;                 assign ID_S_4f622098_66cde942_E[41]  =  6'd53;                 assign ID_S_4f622098_66cde942_E[42]  =  6'd59;                 assign ID_S_4f622098_66cde942_E[43]  =  6'd60;                 assign ID_S_4f622098_66cde942_E[44]  =  6'd30;                 assign ID_S_4f622098_66cde942_E[45]  =  6'd15;                 assign ID_S_4f622098_66cde942_E[46]  =  6'd38;                 assign ID_S_4f622098_66cde942_E[47]  =  6'd19;             end               4'd7:             begin                  assign ID_S_4f622098_66cde942_E[0 ]  =  7'd1;                 assign ID_S_4f622098_66cde942_E[1 ]  =  7'd68;                 assign ID_S_4f622098_66cde942_E[2 ]  =  7'd34;                 assign ID_S_4f622098_66cde942_E[3 ]  =  7'd17;                  assign ID_S_4f622098_66cde942_E[4 ]  =  7'd76;                 assign ID_S_4f622098_66cde942_E[5 ]  =  7'd38;                 assign ID_S_4f622098_66cde942_E[6 ]  =  7'd19;                 assign ID_S_4f622098_66cde942_E[7 ]  =  7'd77;                  assign ID_S_4f622098_66cde942_E[8 ]  =  7'd98;                 assign ID_S_4f622098_66cde942_E[9 ]  =  7'd49;                 assign ID_S_4f622098_66cde942_E[10]  =  7'd92;                 assign ID_S_4f622098_66cde942_E[11]  =  7'd46;                  assign ID_S_4f622098_66cde942_E[12]  =  7'd23;                 assign ID_S_4f622098_66cde942_E[13]  =  7'd79;                 assign ID_S_4f622098_66cde942_E[14]  =  7'd99;                 assign ID_S_4f622098_66cde942_E[15]  =  7'd117;                                                          assign ID_S_4f622098_66cde942_E[16]  =  7'd126;                                 assign ID_S_4f622098_66cde942_E[17]  =  7'd63;                 assign ID_S_4f622098_66cde942_E[18]  =  7'd91;                 assign ID_S_4f622098_66cde942_E[19]  =  7'd105;                 assign ID_S_4f622098_66cde942_E[20]  =  7'd112;                 assign ID_S_4f622098_66cde942_E[21]  =  7'd56;                 assign ID_S_4f622098_66cde942_E[22]  =  7'd28;                 assign ID_S_4f622098_66cde942_E[23]  =  7'd14;                 assign ID_S_4f622098_66cde942_E[24]  =  7'd7;                 assign ID_S_4f622098_66cde942_E[25]  =  7'd71;                 assign ID_S_4f622098_66cde942_E[26]  =  7'd103;                 assign ID_S_4f622098_66cde942_E[27]  =  7'd119;                 assign ID_S_4f622098_66cde942_E[28]  =  7'd127;                 assign ID_S_4f622098_66cde942_E[29]  =  7'd123;                 assign ID_S_4f622098_66cde942_E[30]  =  7'd121;                 assign ID_S_4f622098_66cde942_E[31]  =  7'd120;                                                          assign ID_S_4f622098_66cde942_E[32]  =  7'd60;                 assign ID_S_4f622098_66cde942_E[33]  =  7'd30;                 assign ID_S_4f622098_66cde942_E[34]  =  7'd15;                 assign ID_S_4f622098_66cde942_E[35]  =  7'd67;                 assign ID_S_4f622098_66cde942_E[36]  =  7'd101;                 assign ID_S_4f622098_66cde942_E[37]  =  7'd118;                 assign ID_S_4f622098_66cde942_E[38]  =  7'd59;                 assign ID_S_4f622098_66cde942_E[39]  =  7'd89;                 assign ID_S_4f622098_66cde942_E[40]  =  7'd104;                 assign ID_S_4f622098_66cde942_E[41]  =  7'd52;                 assign ID_S_4f622098_66cde942_E[42]  =  7'd26;                 assign ID_S_4f622098_66cde942_E[43]  =  7'd13;                 assign ID_S_4f622098_66cde942_E[44]  =  7'd66;                 assign ID_S_4f622098_66cde942_E[45]  =  7'd33;                 assign ID_S_4f622098_66cde942_E[46]  =  7'd84;                 assign ID_S_4f622098_66cde942_E[47]  =  7'd42;             end                  4'd8:             begin                  assign ID_S_4f622098_66cde942_E[0 ]  =  8'd1  ;                 assign ID_S_4f622098_66cde942_E[1 ]  =  8'd142;                 assign ID_S_4f622098_66cde942_E[2 ]  =  8'd71 ;                 assign ID_S_4f622098_66cde942_E[3 ]  =  8'd173;                  assign ID_S_4f622098_66cde942_E[4 ]  =  8'd216;                 assign ID_S_4f622098_66cde942_E[5 ]  =  8'd108;                 assign ID_S_4f622098_66cde942_E[6 ]  =  8'd54 ;                 assign ID_S_4f622098_66cde942_E[7 ]  =  8'd27 ;                  assign ID_S_4f622098_66cde942_E[8 ]  =  8'd131;                 assign ID_S_4f622098_66cde942_E[9 ]  =  8'd207;                 assign ID_S_4f622098_66cde942_E[10]  =  8'd233;                 assign ID_S_4f622098_66cde942_E[11]  =  8'd250;                  assign ID_S_4f622098_66cde942_E[12]  =  8'd125;                 assign ID_S_4f622098_66cde942_E[13]  =  8'd176;                 assign ID_S_4f622098_66cde942_E[14]  =  8'd88;                 assign ID_S_4f622098_66cde942_E[15]  =  8'd44;                                    assign ID_S_4f622098_66cde942_E[16]  =  8'd22;                                 assign ID_S_4f622098_66cde942_E[17]  =  8'd11;                 assign ID_S_4f622098_66cde942_E[18]  =  8'd139;                 assign ID_S_4f622098_66cde942_E[19]  =  8'd203;                 assign ID_S_4f622098_66cde942_E[20]  =  8'd235;                 assign ID_S_4f622098_66cde942_E[21]  =  8'd251;                 assign ID_S_4f622098_66cde942_E[22]  =  8'd243;                 assign ID_S_4f622098_66cde942_E[23]  =  8'd247;                 assign ID_S_4f622098_66cde942_E[24]  =  8'd245;                 assign ID_S_4f622098_66cde942_E[25]  =  8'd244;                 assign ID_S_4f622098_66cde942_E[26]  =  8'd122;                 assign ID_S_4f622098_66cde942_E[27]  =  8'd61;                 assign ID_S_4f622098_66cde942_E[28]  =  8'd144;                 assign ID_S_4f622098_66cde942_E[29]  =  8'd72;                 assign ID_S_4f622098_66cde942_E[30]  =  8'd36;                 assign ID_S_4f622098_66cde942_E[31]  =  8'd18;                                   assign ID_S_4f622098_66cde942_E[32]  =  8'd9;                 assign ID_S_4f622098_66cde942_E[33]  =  8'd138;                 assign ID_S_4f622098_66cde942_E[34]  =  8'd69;                 assign ID_S_4f622098_66cde942_E[35]  =  8'd172;                 assign ID_S_4f622098_66cde942_E[36]  =  8'd86;                 assign ID_S_4f622098_66cde942_E[37]  =  8'd43;                 assign ID_S_4f622098_66cde942_E[38]  =  8'd155;                 assign ID_S_4f622098_66cde942_E[39]  =  8'd195;                 assign ID_S_4f622098_66cde942_E[40]  =  8'd239;                 assign ID_S_4f622098_66cde942_E[41]  =  8'd249;                 assign ID_S_4f622098_66cde942_E[42]  =  8'd242;                 assign ID_S_4f622098_66cde942_E[43]  =  8'd121;                 assign ID_S_4f622098_66cde942_E[44]  =  8'd178;                 assign ID_S_4f622098_66cde942_E[45]  =  8'd89;                 assign ID_S_4f622098_66cde942_E[46]  =  8'd162;                 assign ID_S_4f622098_66cde942_E[47]  =  8'd81;             end                     endcase endgenerate          generate     for(ID_S_6227abb2_151191de_E = 0;ID_S_6227abb2_151191de_E <= T_NUM   ;ID_S_6227abb2_151191de_E = ID_S_6227abb2_151191de_E + 1)     begin         case({SYM_BW})             {4'd3}:             begin:ID_S_746774b4_578be916_E                 gf8mul_dec ID_S_636bb82b_1ce12ccd_E   ( ID_S_1cc09e76_634c0c8c_E[ID_S_6227abb2_151191de_E ] ,  ID_S_4f622098_66cde942_E[ID_S_6227abb2_151191de_E]  , ID_S_1439373b_2f1ff4ba_E[ID_S_6227abb2_151191de_E ]);                      end                                                                                    {4'd4}:                                                                                begin:ID_S_4f056043_2154e774_E                                                                         gf16mul_dec ID_S_636bb82b_1ce12ccd_E  ( ID_S_1cc09e76_634c0c8c_E[ID_S_6227abb2_151191de_E ] ,  ID_S_4f622098_66cde942_E[ID_S_6227abb2_151191de_E]  , ID_S_1439373b_2f1ff4ba_E[ID_S_6227abb2_151191de_E ]);                      end                                                                                    {4'd5}:                                                                                begin:ID_S_528be81_2fdc0cc2_E                                                                         gf32mul_dec ID_S_636bb82b_1ce12ccd_E  ( ID_S_1cc09e76_634c0c8c_E[ID_S_6227abb2_151191de_E ] ,  ID_S_4f622098_66cde942_E[ID_S_6227abb2_151191de_E]  , ID_S_1439373b_2f1ff4ba_E[ID_S_6227abb2_151191de_E ]);                      end                                                                                    {4'd6}:                                                                                begin:ID_S_7a4153e6_3d475d01_E                                                                         gf64mul_dec ID_S_636bb82b_1ce12ccd_E  ( ID_S_1cc09e76_634c0c8c_E[ID_S_6227abb2_151191de_E ] ,  ID_S_4f622098_66cde942_E[ID_S_6227abb2_151191de_E]  , ID_S_1439373b_2f1ff4ba_E[ID_S_6227abb2_151191de_E ]);                      end                                                                                    {4'd7}:                                                                                begin:ID_S_72795317_48c1aab1_E                                                                        gf128mul_dec ID_S_636bb82b_1ce12ccd_E ( ID_S_1cc09e76_634c0c8c_E[ID_S_6227abb2_151191de_E ] ,  ID_S_4f622098_66cde942_E[ID_S_6227abb2_151191de_E]  , ID_S_1439373b_2f1ff4ba_E[ID_S_6227abb2_151191de_E ]);                      end                                                                                                                                                                           {4'd8}:                                                                                begin:ID_S_1afcd9b9_23d4718d_E                                                                        gf256mul_dec ID_S_636bb82b_1ce12ccd_E ( ID_S_1cc09e76_634c0c8c_E[ID_S_6227abb2_151191de_E ] ,  ID_S_4f622098_66cde942_E[ID_S_6227abb2_151191de_E]  , ID_S_1439373b_2f1ff4ba_E[ID_S_6227abb2_151191de_E ]);                     end         endcase                   end endgenerate  generate     for(ID_S_6227abb2_151191de_E = 0;ID_S_6227abb2_151191de_E < T_NUM   ;ID_S_6227abb2_151191de_E = ID_S_6227abb2_151191de_E + 1)     begin         case({SYM_BW})             {4'd3}:             begin:ID_S_746774b5_578be915_E                 gf8mul_dec ID_S_637dd0ac_1c136950_E   ( ID_S_34d46d67_7fcdf326_E[ID_S_6227abb2_151191de_E] ,  ID_S_4f622098_66cde942_E[2*T_NUM + ID_S_6227abb2_151191de_E] , ID_S_763fe6b_156a0a07_E[ID_S_6227abb2_151191de_E ]);             end                                                              {4'd4}:                                                          begin:ID_S_4f056044_2154e777_E                                                   gf16mul_dec ID_S_637dd0ac_1c136950_E  ( ID_S_34d46d67_7fcdf326_E[ID_S_6227abb2_151191de_E] ,  ID_S_4f622098_66cde942_E[2*T_NUM + ID_S_6227abb2_151191de_E] , ID_S_763fe6b_156a0a07_E[ID_S_6227abb2_151191de_E ]);             end                                                              {4'd5}:                                                          begin:ID_S_528be82_2fdc0cc1_E                                                   gf32mul_dec ID_S_637dd0ac_1c136950_E  ( ID_S_34d46d67_7fcdf326_E[ID_S_6227abb2_151191de_E] ,  ID_S_4f622098_66cde942_E[2*T_NUM + ID_S_6227abb2_151191de_E] , ID_S_763fe6b_156a0a07_E[ID_S_6227abb2_151191de_E ]);             end                                                              {4'd6}:                                                          begin:ID_S_7a4153e7_3d475d02_E                                                   gf64mul_dec ID_S_637dd0ac_1c136950_E  ( ID_S_34d46d67_7fcdf326_E[ID_S_6227abb2_151191de_E] ,  ID_S_4f622098_66cde942_E[2*T_NUM + ID_S_6227abb2_151191de_E] , ID_S_763fe6b_156a0a07_E[ID_S_6227abb2_151191de_E ]);             end                                                              {4'd7}:                                                          begin:ID_S_72795318_48c1aab2_E                                                  gf128mul_dec ID_S_637dd0ac_1c136950_E ( ID_S_34d46d67_7fcdf326_E[ID_S_6227abb2_151191de_E] ,  ID_S_4f622098_66cde942_E[2*T_NUM + ID_S_6227abb2_151191de_E] , ID_S_763fe6b_156a0a07_E[ID_S_6227abb2_151191de_E ]);             end                                                                                                                               {4'd8}:                                                          begin:ID_S_1afcd9ba_23d4718e_E                                                  gf256mul_dec ID_S_637dd0ac_1c136950_E ( ID_S_34d46d67_7fcdf326_E[ID_S_6227abb2_151191de_E] ,  ID_S_4f622098_66cde942_E[2*T_NUM + ID_S_6227abb2_151191de_E] , ID_S_763fe6b_156a0a07_E[ID_S_6227abb2_151191de_E ]);             end         endcase                   end endgenerate   generate     for(ID_S_6227abb2_151191de_E = 0;ID_S_6227abb2_151191de_E < T_NUM   ;ID_S_6227abb2_151191de_E = ID_S_6227abb2_151191de_E + 1)     begin         always @(posedge clk or negedge rst_n)         if (!rst_n)         begin           ID_S_34d46d67_7fcdf326_E[ID_S_6227abb2_151191de_E] <= 0;         end         else if (start)         begin           ID_S_34d46d67_7fcdf326_E[ID_S_6227abb2_151191de_E]       <= 8'd1;         end         else if (ID_S_651d5efd_799ab730_E)         begin           ID_S_34d46d67_7fcdf326_E[ID_S_6227abb2_151191de_E]       <= ID_S_763fe6b_156a0a07_E[ID_S_6227abb2_151191de_E]      ;          end         else         begin           ID_S_34d46d67_7fcdf326_E[ID_S_6227abb2_151191de_E]       <= 0;          end             end endgenerate    generate     for(ID_S_6227abb2_151191de_E = 0;ID_S_6227abb2_151191de_E <= T_NUM   ;ID_S_6227abb2_151191de_E = ID_S_6227abb2_151191de_E + 1)     begin         always @(posedge clk or negedge rst_n)         if (!rst_n)         begin           ID_S_1cc09e76_634c0c8c_E[ID_S_6227abb2_151191de_E] <= 0;         end         else if (start)         begin           ID_S_1cc09e76_634c0c8c_E[ID_S_6227abb2_151191de_E]       <= 8'd1;         end         else if (ID_S_651d5efd_799ab730_E)         begin           ID_S_1cc09e76_634c0c8c_E[ID_S_6227abb2_151191de_E]       <= ID_S_1439373b_2f1ff4ba_E[ID_S_6227abb2_151191de_E]      ;         end         else         begin           ID_S_1cc09e76_634c0c8c_E[ID_S_6227abb2_151191de_E]       <= 0      ;         end             end endgenerate   wire [SYM_BW-1:0] ID_S_630efec2_48bceb62_E[ID_S_b8824c0_7ead0f40_E - 1:0]; wire [SYM_BW-1:0] ID_S_4485e2ac_30899592_E[T_NUM - 1:0];  generate     for(ID_S_6227abb2_151191de_E = 0;ID_S_6227abb2_151191de_E < T_NUM   ;ID_S_6227abb2_151191de_E = ID_S_6227abb2_151191de_E + 1)     begin         case({SYM_BW})             {4'd3}:             begin:ID_S_746774b6_578be914_E                 gf8mul_dec ID_S_ea35e67_7effe83_E  ( ID_S_34d46d67_7fcdf326_E[ID_S_6227abb2_151191de_E] ,  ID_S_69e010d1_7dab0633_E[ID_S_6227abb2_151191de_E], ID_S_4485e2ac_30899592_E[ID_S_6227abb2_151191de_E]);                             end                                                          {4'd4}:                                                      begin:ID_S_4f056045_2154e776_E                                               gf16mul_dec ID_S_ea35e67_7effe83_E ( ID_S_34d46d67_7fcdf326_E[ID_S_6227abb2_151191de_E] ,  ID_S_69e010d1_7dab0633_E[ID_S_6227abb2_151191de_E], ID_S_4485e2ac_30899592_E[ID_S_6227abb2_151191de_E]);                             end                                                          {4'd5}:                                                      begin:ID_S_528be83_2fdc0cc0_E                                               gf32mul_dec ID_S_ea35e67_7effe83_E ( ID_S_34d46d67_7fcdf326_E[ID_S_6227abb2_151191de_E] ,  ID_S_69e010d1_7dab0633_E[ID_S_6227abb2_151191de_E], ID_S_4485e2ac_30899592_E[ID_S_6227abb2_151191de_E]);                             end                                                          {4'd6}:                                                      begin:ID_S_7a4153e8_3d475d03_E                                               gf64mul_dec ID_S_ea35e67_7effe83_E ( ID_S_34d46d67_7fcdf326_E[ID_S_6227abb2_151191de_E] ,  ID_S_69e010d1_7dab0633_E[ID_S_6227abb2_151191de_E], ID_S_4485e2ac_30899592_E[ID_S_6227abb2_151191de_E]);                             end                                                          {4'd7}:                                                      begin:ID_S_72795319_48c1aab3_E                                              gf128mul_dec ID_S_ea35e67_7effe83_E( ID_S_34d46d67_7fcdf326_E[ID_S_6227abb2_151191de_E] ,  ID_S_69e010d1_7dab0633_E[ID_S_6227abb2_151191de_E], ID_S_4485e2ac_30899592_E[ID_S_6227abb2_151191de_E]);                             end                                                                                                                       {4'd8}:                                                      begin:ID_S_1afcd9bb_23d4718f_E                                              gf256mul_dec ID_S_ea35e67_7effe83_E( ID_S_34d46d67_7fcdf326_E[ID_S_6227abb2_151191de_E] ,  ID_S_69e010d1_7dab0633_E[ID_S_6227abb2_151191de_E], ID_S_4485e2ac_30899592_E[ID_S_6227abb2_151191de_E]);                             end         endcase                   end endgenerate  generate     for(ID_S_6227abb2_151191de_E = 1;ID_S_6227abb2_151191de_E <= T_NUM   ;ID_S_6227abb2_151191de_E = ID_S_6227abb2_151191de_E + 2)     begin         case({SYM_BW})             {4'd3}:             begin:ID_S_746774b7_578be913_E                 gf8mul_dec ID_S_ea35e46_7efc684_E  (ID_S_1cc09e76_634c0c8c_E[ID_S_6227abb2_151191de_E] , ID_S_678291e7_5121332d_E[ID_S_6227abb2_151191de_E], ID_S_630efec2_48bceb62_E[(ID_S_6227abb2_151191de_E-1)/2]);             end                                                       {4'd4}:                                                   begin:ID_S_4f056046_2154e771_E                                            gf16mul_dec ID_S_ea35e46_7efc684_E (ID_S_1cc09e76_634c0c8c_E[ID_S_6227abb2_151191de_E] , ID_S_678291e7_5121332d_E[ID_S_6227abb2_151191de_E], ID_S_630efec2_48bceb62_E[(ID_S_6227abb2_151191de_E-1)/2]);             end                                                       {4'd5}:                                                   begin:ID_S_528be84_2fdc0cc7_E                                            gf32mul_dec ID_S_ea35e46_7efc684_E (ID_S_1cc09e76_634c0c8c_E[ID_S_6227abb2_151191de_E] , ID_S_678291e7_5121332d_E[ID_S_6227abb2_151191de_E], ID_S_630efec2_48bceb62_E[(ID_S_6227abb2_151191de_E-1)/2]);             end                                                       {4'd6}:                                                   begin:ID_S_7a4153e9_3d475d04_E                                            gf64mul_dec ID_S_ea35e46_7efc684_E (ID_S_1cc09e76_634c0c8c_E[ID_S_6227abb2_151191de_E] , ID_S_678291e7_5121332d_E[ID_S_6227abb2_151191de_E], ID_S_630efec2_48bceb62_E[(ID_S_6227abb2_151191de_E-1)/2]);             end                                                       {4'd7}:                                                   begin:ID_S_7279531a_48c1aab4_E                                           gf128mul_dec ID_S_ea35e46_7efc684_E(ID_S_1cc09e76_634c0c8c_E[ID_S_6227abb2_151191de_E] , ID_S_678291e7_5121332d_E[ID_S_6227abb2_151191de_E], ID_S_630efec2_48bceb62_E[(ID_S_6227abb2_151191de_E-1)/2]);             end                                                                                                                 {4'd8}:                                                   begin:ID_S_1afcd9bc_23d47188_E                                           gf256mul_dec ID_S_ea35e46_7efc684_E(ID_S_1cc09e76_634c0c8c_E[ID_S_6227abb2_151191de_E] , ID_S_678291e7_5121332d_E[ID_S_6227abb2_151191de_E], ID_S_630efec2_48bceb62_E[(ID_S_6227abb2_151191de_E-1)/2]);             end         endcase                   end endgenerate        reg [SYM_BW-1:0] ID_S_57d4d0a8_25cef536_E; reg [SYM_BW-1:0] ID_S_69e010e3_7dab0621_E;  wire [SYM_BW-1:0] ID_S_204ba75e_59c45ac1_E; wire [SYM_BW-1:0] ID_S_6227e259_156d64f1_E;  generate     case({T_NUM})         {
`R_BW'd1}:

        begin:ID_S_1c3375e2_144f0e9e_E             assign ID_S_204ba75e_59c45ac1_E = ID_S_630efec2_48bceb62_E[0]  ;             assign ID_S_6227e259_156d64f1_E  = ID_S_4485e2ac_30899592_E[0]  ;         end             {
`R_BW'd2}:

        begin:ID_S_1c3375e3_144f0e9d_E             assign ID_S_204ba75e_59c45ac1_E = ID_S_630efec2_48bceb62_E[0]  ;             assign ID_S_6227e259_156d64f1_E  = ID_S_4485e2ac_30899592_E[0] ^ ID_S_4485e2ac_30899592_E[1] ;         end         {
`R_BW'd4}:

        begin:ID_S_1c3375e5_144f0e9b_E             assign ID_S_204ba75e_59c45ac1_E = ID_S_630efec2_48bceb62_E[0] ^ ID_S_630efec2_48bceb62_E[1] ;             assign ID_S_6227e259_156d64f1_E  = ID_S_4485e2ac_30899592_E[0] ^ ID_S_4485e2ac_30899592_E[1] ^ ID_S_4485e2ac_30899592_E[2] ^ ID_S_4485e2ac_30899592_E[3] ;         end                           {
`R_BW'd8}:

        begin:ID_S_1c3375e9_144f0e97_E             assign ID_S_204ba75e_59c45ac1_E = ID_S_630efec2_48bceb62_E[0] ^ ID_S_630efec2_48bceb62_E[1] ^ ID_S_630efec2_48bceb62_E[2] ^ ID_S_630efec2_48bceb62_E[3];             assign ID_S_6227e259_156d64f1_E  = ID_S_4485e2ac_30899592_E[0] ^ ID_S_4485e2ac_30899592_E[1] ^ ID_S_4485e2ac_30899592_E[2] ^ ID_S_4485e2ac_30899592_E[3] ^ ID_S_4485e2ac_30899592_E[4] ^ ID_S_4485e2ac_30899592_E[5] ^ ID_S_4485e2ac_30899592_E[6] ^ ID_S_4485e2ac_30899592_E[7];         end         {
`R_BW'd16}:

        begin:ID_S_22a23258_13667923_E             assign ID_S_204ba75e_59c45ac1_E = ID_S_630efec2_48bceb62_E[0] ^ ID_S_630efec2_48bceb62_E[1] ^ ID_S_630efec2_48bceb62_E[2] ^ ID_S_630efec2_48bceb62_E[3] ^ ID_S_630efec2_48bceb62_E[4] ^ ID_S_630efec2_48bceb62_E[5] ^ ID_S_630efec2_48bceb62_E[6] ^ ID_S_630efec2_48bceb62_E[7];             assign ID_S_6227e259_156d64f1_E  = ID_S_4485e2ac_30899592_E[0] ^ ID_S_4485e2ac_30899592_E[1] ^ ID_S_4485e2ac_30899592_E[2] ^ ID_S_4485e2ac_30899592_E[3] ^ ID_S_4485e2ac_30899592_E[4] ^ ID_S_4485e2ac_30899592_E[5] ^ ID_S_4485e2ac_30899592_E[6] ^ ID_S_4485e2ac_30899592_E[7] ^ ID_S_4485e2ac_30899592_E[8] ^ ID_S_4485e2ac_30899592_E[9] ^ ID_S_4485e2ac_30899592_E[10] ^ ID_S_4485e2ac_30899592_E[11] ^ ID_S_4485e2ac_30899592_E[12] ^ ID_S_4485e2ac_30899592_E[13] ^ ID_S_4485e2ac_30899592_E[14] ^ ID_S_4485e2ac_30899592_E[15];         end             endcase endgenerate     always @(posedge clk or negedge rst_n) if (!rst_n) begin     ID_S_57d4d0a8_25cef536_E <= 8'd0;     ID_S_69e010e3_7dab0621_E  <= 8'd0;   end else if (start) begin     ID_S_57d4d0a8_25cef536_E <= 8'd0;     ID_S_69e010e3_7dab0621_E  <= 8'd0;      end else if (ID_S_651d5efd_799ab730_E) begin     ID_S_57d4d0a8_25cef536_E <= ID_S_204ba75e_59c45ac1_E;     ID_S_69e010e3_7dab0621_E  <= ID_S_6227e259_156d64f1_E ; end      wire [SYM_BW-1:0] ID_S_61d2c9f4_4cdb9c10_E;       reg [SYM_BW-1:0]  ID_S_857c936_48fbcfab_E; reg [SYM_BW-1:0]  ID_S_1350f028_6b3eb61b_E; always @(posedge clk or negedge rst_n) if (!rst_n) begin     ID_S_857c936_48fbcfab_E  <= 8'd0; end else  begin     ID_S_857c936_48fbcfab_E  <= N_NUM + 1 - ID_S_651d5efd_799ab730_E ;   end  always @(posedge clk or negedge rst_n) if (!rst_n) begin     ID_S_1350f028_6b3eb61b_E  <= 8'd0; end else  begin     ID_S_1350f028_6b3eb61b_E  <= {{(8-SYM_BW){1'b0}},{SYM_BW{1'b1}}} + 8'd1 - ID_S_651d5efd_799ab730_E ;   end   wire [SYM_BW-1:0] ID_S_77b0927b_625887db_E; wire [SYM_BW-1:0] ID_S_4129a3aa_30f01dd2_E; wire [SYM_BW-1:0] ID_S_15169203_bbc8e76_E;  generate         case({SYM_BW})         {4'd3}:         begin:gf8inv             gf8inv ID_S_7e3fbf2b_1b2ada90_E( ID_S_57d4d0a8_25cef536_E, ID_S_61d2c9f4_4cdb9c10_E);               idx2gf8 ID_S_5fe9a495_74a16f65_E( ID_S_1350f028_6b3eb61b_E, ID_S_77b0927b_625887db_E);             gf8mul_dec ID_S_ea35e88_7eff682_E(ID_S_69e010e3_7dab0621_E, ID_S_61d2c9f4_4cdb9c10_E, ID_S_4129a3aa_30f01dd2_E);             gf8mul_dec ID_S_ea35ea9_7efee81_E(ID_S_4129a3aa_30f01dd2_E, ID_S_77b0927b_625887db_E, ID_S_15169203_bbc8e76_E);         end         {4'd4}:         begin:gf16inv             gf16inv ID_S_7e3fbf2b_1b2ada90_E( ID_S_57d4d0a8_25cef536_E, ID_S_61d2c9f4_4cdb9c10_E);               idx2gf16 ID_S_5fe9a495_74a16f65_E( ID_S_1350f028_6b3eb61b_E, ID_S_77b0927b_625887db_E);             gf16mul_dec ID_S_ea35e88_7eff682_E(ID_S_69e010e3_7dab0621_E, ID_S_61d2c9f4_4cdb9c10_E, ID_S_4129a3aa_30f01dd2_E);             gf16mul_dec ID_S_ea35ea9_7efee81_E(ID_S_4129a3aa_30f01dd2_E, ID_S_77b0927b_625887db_E, ID_S_15169203_bbc8e76_E);         end         {4'd5}:         begin:gf32inv             gf32inv ID_S_7e3fbf2b_1b2ada90_E( ID_S_57d4d0a8_25cef536_E, ID_S_61d2c9f4_4cdb9c10_E);               idx2gf32 ID_S_5fe9a495_74a16f65_E( ID_S_1350f028_6b3eb61b_E, ID_S_77b0927b_625887db_E);             gf32mul_dec ID_S_ea35e88_7eff682_E(ID_S_69e010e3_7dab0621_E, ID_S_61d2c9f4_4cdb9c10_E, ID_S_4129a3aa_30f01dd2_E);             gf32mul_dec ID_S_ea35ea9_7efee81_E(ID_S_4129a3aa_30f01dd2_E, ID_S_77b0927b_625887db_E, ID_S_15169203_bbc8e76_E);         end         {4'd6}:         begin:gf64inv             gf64inv ID_S_7e3fbf2b_1b2ada90_E( ID_S_57d4d0a8_25cef536_E, ID_S_61d2c9f4_4cdb9c10_E);               idx2gf64 ID_S_5fe9a495_74a16f65_E( ID_S_1350f028_6b3eb61b_E, ID_S_77b0927b_625887db_E);             gf64mul_dec ID_S_ea35e88_7eff682_E(ID_S_69e010e3_7dab0621_E, ID_S_61d2c9f4_4cdb9c10_E, ID_S_4129a3aa_30f01dd2_E);             gf64mul_dec ID_S_ea35ea9_7efee81_E(ID_S_4129a3aa_30f01dd2_E, ID_S_77b0927b_625887db_E, ID_S_15169203_bbc8e76_E);         end         {4'd7}:         begin:gf128inv             gf128inv ID_S_7e3fbf2b_1b2ada90_E( ID_S_57d4d0a8_25cef536_E, ID_S_61d2c9f4_4cdb9c10_E);               idx2gf128 ID_S_5fe9a495_74a16f65_E( ID_S_1350f028_6b3eb61b_E, ID_S_77b0927b_625887db_E);             gf128mul_dec ID_S_ea35e88_7eff682_E(ID_S_69e010e3_7dab0621_E, ID_S_61d2c9f4_4cdb9c10_E, ID_S_4129a3aa_30f01dd2_E);             gf128mul_dec ID_S_ea35ea9_7efee81_E(ID_S_4129a3aa_30f01dd2_E, ID_S_77b0927b_625887db_E, ID_S_15169203_bbc8e76_E);         end                   {4'd8}:         begin:gf256inv             gf256inv ID_S_7b616a10_1cb5d2e3_E( ID_S_57d4d0a8_25cef536_E, ID_S_61d2c9f4_4cdb9c10_E);               idx2gf256 ID_S_e50b5a_40011093_E( ID_S_1350f028_6b3eb61b_E, ID_S_77b0927b_625887db_E);             gf256mul_dec ID_S_ea35e88_7eff682_E(ID_S_69e010e3_7dab0621_E, ID_S_61d2c9f4_4cdb9c10_E, ID_S_4129a3aa_30f01dd2_E);             gf256mul_dec ID_S_ea35ea9_7efee81_E(ID_S_4129a3aa_30f01dd2_E, ID_S_77b0927b_625887db_E, ID_S_15169203_bbc8e76_E);                      end     endcase     endgenerate  generate     for(ID_S_6227abb2_151191de_E = 0;ID_S_6227abb2_151191de_E < T_NUM  ;ID_S_6227abb2_151191de_E = ID_S_6227abb2_151191de_E + 1)     begin         always @(posedge clk or negedge rst_n)         if (!rst_n)         begin             err_val[(ID_S_6227abb2_151191de_E+1) *SYM_BW - 1:ID_S_6227abb2_151191de_E *SYM_BW] <= 8'd0;             err_loc_out[(ID_S_6227abb2_151191de_E+1) *SYM_BW - 1:ID_S_6227abb2_151191de_E *SYM_BW] <= 8'd0;         end else if (start) begin             err_val[(ID_S_6227abb2_151191de_E+1) *SYM_BW - 1:ID_S_6227abb2_151191de_E *SYM_BW] <= 8'd0;             err_loc_out[(ID_S_6227abb2_151191de_E+1) *SYM_BW - 1:ID_S_6227abb2_151191de_E *SYM_BW] <= 8'd0;         end else if (ID_S_857c936_48fbcfab_E) begin             case(ID_S_857c936_48fbcfab_E)                 ID_S_496ff42e_ba097b9_E[ID_S_6227abb2_151191de_E]:                       begin                          err_val[(ID_S_6227abb2_151191de_E+1) *SYM_BW - 1: ID_S_6227abb2_151191de_E*SYM_BW] <=  ID_S_15169203_bbc8e76_E;                             err_loc_out[(ID_S_6227abb2_151191de_E+1) *SYM_BW - 1: ID_S_6227abb2_151191de_E*SYM_BW]  <= ID_S_857c936_48fbcfab_E;                      end                 default:;             endcase         end else              ;             end endgenerate    reg ID_S_69599382_7da7a65d_E; always @(posedge clk or negedge rst_n) if (!rst_n)     ID_S_69599382_7da7a65d_E <= 0; else if (ID_S_651d5efd_799ab730_E == N_NUM)     ID_S_69599382_7da7a65d_E <= 1; else     ID_S_69599382_7da7a65d_E <= 0;  always @(posedge clk or negedge rst_n) if (!rst_n)     done <= 0; else     done <= ID_S_69599382_7da7a65d_E;      endmodule  