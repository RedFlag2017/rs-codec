`timescale 1ns/100ps
module gf32mul(
    input       [4:0] a,
    input       [4:0] b,
    output  reg [4:0] z
);
always @(*)
begin
    case (b)
        5'd1:
            begin
                z[0] = a[0];
                z[1] = a[1];
                z[2] = a[2];
                z[3] = a[3];
                z[4] = a[4];
            end
        5'd2:
            begin
                z[0] = a[4];
                z[1] = a[0];
                z[2] = a[1] ^ a[4];
                z[3] = a[2];
                z[4] = a[3];
            end
        5'd3:
            begin
                z[0] = a[0] ^ a[4];
                z[1] = a[0] ^ a[1];
                z[2] = a[1] ^ a[2] ^ a[4];
                z[3] = a[2] ^ a[3];
                z[4] = a[3] ^ a[4];
            end
        5'd5:
            begin
                z[0] = a[0] ^ a[3];
                z[1] = a[1] ^ a[4];
                z[2] = a[0] ^ a[2] ^ a[3];
                z[3] = a[1] ^ a[3] ^ a[4];
                z[4] = a[2] ^ a[4];
            end
        5'd6:
            begin
                z[0] = a[3] ^ a[4];
                z[1] = a[0] ^ a[4];
                z[2] = a[0] ^ a[1] ^ a[3] ^ a[4];
                z[3] = a[1] ^ a[2] ^ a[4];
                z[4] = a[2] ^ a[3];
            end
        5'd8:
            begin
                z[0] = a[2];
                z[1] = a[3];
                z[2] = a[2] ^ a[4];
                z[3] = a[0] ^ a[3];
                z[4] = a[1] ^ a[4];
            end
        5'd9:
            begin
                z[0] = a[0] ^ a[2];
                z[1] = a[1] ^ a[3];
                z[2] = a[4];
                z[3] = a[0];
                z[4] = a[1];
            end
        5'd13:
            begin
                z[0] = a[0] ^ a[2] ^ a[3];
                z[1] = a[1] ^ a[3] ^ a[4];
                z[2] = a[0] ^ a[3] ^ a[4];
                z[3] = a[0] ^ a[1] ^ a[4];
                z[4] = a[1] ^ a[2];
            end
        5'd14:
            begin
                z[0] = a[2] ^ a[3] ^ a[4];
                z[1] = a[0] ^ a[3] ^ a[4];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[3];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
                z[4] = a[1] ^ a[2] ^ a[3] ^ a[4];
            end
        5'd15:
            begin
                z[0] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[1] = a[0] ^ a[1] ^ a[3] ^ a[4];
                z[2] = a[0] ^ a[1] ^ a[3];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[4];
                z[4] = a[1] ^ a[2] ^ a[3];
            end
        5'd16:
            begin
                z[0] = a[1] ^ a[4];
                z[1] = a[2];
                z[2] = a[1] ^ a[3] ^ a[4];
                z[3] = a[2] ^ a[4];
                z[4] = a[0] ^ a[3];
            end
        5'd17:
            begin
                z[0] = a[0] ^ a[1] ^ a[4];
                z[1] = a[1] ^ a[2];
                z[2] = a[1] ^ a[2] ^ a[3] ^ a[4];
                z[3] = a[2] ^ a[3] ^ a[4];
                z[4] = a[0] ^ a[3] ^ a[4];
            end
        5'd18:
            begin
                z[0] = a[1];
                z[1] = a[0] ^ a[2];
                z[2] = a[3];
                z[3] = a[4];
                z[4] = a[0];
            end
        5'd20:
            begin
                z[0] = a[1] ^ a[3] ^ a[4];
                z[1] = a[2] ^ a[4];
                z[2] = a[0] ^ a[1] ^ a[4];
                z[3] = a[1] ^ a[2];
                z[4] = a[0] ^ a[2] ^ a[3];
            end
        5'd21:
            begin
                z[0] = a[0] ^ a[1] ^ a[3] ^ a[4];
                z[1] = a[1] ^ a[2] ^ a[4];
                z[2] = a[0] ^ a[1] ^ a[2] ^ a[4];
                z[3] = a[1] ^ a[2] ^ a[3];
                z[4] = a[0] ^ a[2] ^ a[3] ^ a[4];
            end
        5'd24:
            begin
                z[0] = a[1] ^ a[2] ^ a[4];
                z[1] = a[2] ^ a[3];
                z[2] = a[1] ^ a[2] ^ a[3];
                z[3] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[4] = a[0] ^ a[1] ^ a[3] ^ a[4];
            end
        5'd25:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[4];
                z[1] = a[1] ^ a[2] ^ a[3];
                z[2] = a[1] ^ a[3];
                z[3] = a[0] ^ a[2] ^ a[4];
                z[4] = a[0] ^ a[1] ^ a[3];
            end
        5'd26:
            begin
                z[0] = a[1] ^ a[2];
                z[1] = a[0] ^ a[2] ^ a[3];
                z[2] = a[2] ^ a[3] ^ a[4];
                z[3] = a[0] ^ a[3] ^ a[4];
                z[4] = a[0] ^ a[1] ^ a[4];
            end
        5'd28:
            begin
                z[0] = a[1] ^ a[2] ^ a[3] ^ a[4];
                z[1] = a[2] ^ a[3] ^ a[4];
                z[2] = a[0] ^ a[1] ^ a[2];
                z[3] = a[0] ^ a[1] ^ a[2] ^ a[3];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
            end
        5'd29:
            begin
                z[0] = a[0] ^ a[1] ^ a[2] ^ a[3] ^ a[4];
                z[1] = a[1] ^ a[2] ^ a[3] ^ a[4];
                z[2] = a[0] ^ a[1];
                z[3] = a[0] ^ a[1] ^ a[2];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[3];
            end
        5'd30:
            begin
                z[0] = a[1] ^ a[2] ^ a[3];
                z[1] = a[0] ^ a[2] ^ a[3] ^ a[4];
                z[2] = a[0] ^ a[2] ^ a[4];
                z[3] = a[0] ^ a[1] ^ a[3];
                z[4] = a[0] ^ a[1] ^ a[2] ^ a[4];
            end
        default:
            begin
                z[0] = 0; 
                z[1] = 0; 
                z[2] = 0; 
                z[3] = 0; 
                z[4] = 0; 
            end
    endcase
end
endmodule
