
`include "smp_if.sv" 
`include "test_collection.sv" 