 
`timescale 1ns/100ps

module rs_lfsr  #( parameter [3:0] SYM_BW = 8, parameter [8-1:0]  N_NUM = 255, parameter [
`R_BW-1:0]  R_NUM = 16

)  (     input clk,     input rst_n,     input din_val,     input din_sop,     input [SYM_BW - 1:0] din,     output reg dout_val,     output reg dout_sop,     output reg dout_eop,     output reg [SYM_BW - 1 :0] dout  );   localparam ID_S_12846e01_7d0ea1dd_E = SYM_BW;   wire [SYM_BW-1:0] ID_S_7f18c66f_6de04cff_E[R_NUM - 1:0]  ;  generate     case({ID_S_12846e01_7d0ea1dd_E,R_NUM})          {4'd3,6'd4}:             begin                  assign ID_S_7f18c66f_6de04cff_E[0]  = 3'd3 ;                 assign ID_S_7f18c66f_6de04cff_E[1]  = 3'd2 ;                 assign ID_S_7f18c66f_6de04cff_E[2]  = 3'd1 ;                 assign ID_S_7f18c66f_6de04cff_E[3]  = 3'd3 ;                      end         {4'd3,6'd3}:             begin                  assign ID_S_7f18c66f_6de04cff_E[0]  = 3'd5 ;                 assign ID_S_7f18c66f_6de04cff_E[1]  = 3'd2 ;                 assign ID_S_7f18c66f_6de04cff_E[2]  = 3'd5 ;             end         {4'd3,6'd2}:             begin                  assign ID_S_7f18c66f_6de04cff_E[0]  = 3'd3 ;                 assign ID_S_7f18c66f_6de04cff_E[1]  = 3'd6 ;             end                                                  {4'd4,6'd2}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 4'd8;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 4'd6;             end          {4'd4,6'd4}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 4'd7;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 4'd8;                 assign ID_S_7f18c66f_6de04cff_E[2 ] = 4'd12;                 assign ID_S_7f18c66f_6de04cff_E[3 ] = 4'd13;             end          {4'd4,6'd8}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 4'd12;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 4'd14;                 assign ID_S_7f18c66f_6de04cff_E[2 ] = 4'd6;                 assign ID_S_7f18c66f_6de04cff_E[3 ] = 4'd13;                 assign ID_S_7f18c66f_6de04cff_E[4 ] = 4'd4;                 assign ID_S_7f18c66f_6de04cff_E[5 ] = 4'd3;                 assign ID_S_7f18c66f_6de04cff_E[6 ] = 4'd4;                 assign ID_S_7f18c66f_6de04cff_E[7 ] = 4'd9;             end                              {4'd5,6'd2}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 5'd8;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 5'd6;             end          {4'd5,6'd4}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 5'd17;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 5'd9;                 assign ID_S_7f18c66f_6de04cff_E[2 ] = 5'd6;                 assign ID_S_7f18c66f_6de04cff_E[3 ] = 5'd30;             end          {4'd5,6'd8}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 5'd5;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 5'd18;                 assign ID_S_7f18c66f_6de04cff_E[2 ] = 5'd26;                 assign ID_S_7f18c66f_6de04cff_E[3 ] = 5'd2;                 assign ID_S_7f18c66f_6de04cff_E[4 ] = 5'd6;                 assign ID_S_7f18c66f_6de04cff_E[5 ] = 5'd15;                 assign ID_S_7f18c66f_6de04cff_E[6 ] = 5'd21;                 assign ID_S_7f18c66f_6de04cff_E[7 ] = 5'd8;             end          {4'd5,6'd16}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 5'd14;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 5'd3;                 assign ID_S_7f18c66f_6de04cff_E[2 ] = 5'd21;                 assign ID_S_7f18c66f_6de04cff_E[3 ] = 5'd15;                 assign ID_S_7f18c66f_6de04cff_E[4 ] = 5'd29;                 assign ID_S_7f18c66f_6de04cff_E[5 ] = 5'd15;                 assign ID_S_7f18c66f_6de04cff_E[6 ] = 5'd16;                 assign ID_S_7f18c66f_6de04cff_E[7 ] = 5'd20;                 assign ID_S_7f18c66f_6de04cff_E[8 ] = 5'd25;                 assign ID_S_7f18c66f_6de04cff_E[9 ] = 5'd24;                 assign ID_S_7f18c66f_6de04cff_E[10] = 5'd2;                 assign ID_S_7f18c66f_6de04cff_E[11] = 5'd8;                 assign ID_S_7f18c66f_6de04cff_E[12] = 5'd13;                 assign ID_S_7f18c66f_6de04cff_E[13] = 5'd1;                 assign ID_S_7f18c66f_6de04cff_E[14] = 5'd28;                 assign ID_S_7f18c66f_6de04cff_E[15] = 5'd15;             end                                   {4'd6,6'd2}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 6'd8;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 6'd6;             end          {4'd6,6'd4}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 6'd48;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 6'd17;                 assign ID_S_7f18c66f_6de04cff_E[2 ] = 6'd29;                 assign ID_S_7f18c66f_6de04cff_E[3 ] = 6'd30;             end          {4'd6,6'd8}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 6'd22;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 6'd6;                 assign ID_S_7f18c66f_6de04cff_E[2 ] = 6'd20;                 assign ID_S_7f18c66f_6de04cff_E[3 ] = 6'd47;                 assign ID_S_7f18c66f_6de04cff_E[4 ] = 6'd48;                 assign ID_S_7f18c66f_6de04cff_E[5 ] = 6'd37;                 assign ID_S_7f18c66f_6de04cff_E[6 ] = 6'd61;                 assign ID_S_7f18c66f_6de04cff_E[7 ] = 6'd55;             end          {4'd6,6'd16}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 6'd48;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 6'd59;                 assign ID_S_7f18c66f_6de04cff_E[2 ] = 6'd38;                 assign ID_S_7f18c66f_6de04cff_E[3 ] = 6'd41;                 assign ID_S_7f18c66f_6de04cff_E[4 ] = 6'd59;                 assign ID_S_7f18c66f_6de04cff_E[5 ] = 6'd5;                 assign ID_S_7f18c66f_6de04cff_E[6 ] = 6'd34;                 assign ID_S_7f18c66f_6de04cff_E[7 ] = 6'd52;                 assign ID_S_7f18c66f_6de04cff_E[8 ] = 6'd27;                 assign ID_S_7f18c66f_6de04cff_E[9 ] = 6'd18;                 assign ID_S_7f18c66f_6de04cff_E[10] = 6'd23;                 assign ID_S_7f18c66f_6de04cff_E[11] = 6'd17;                 assign ID_S_7f18c66f_6de04cff_E[12] = 6'd19;                 assign ID_S_7f18c66f_6de04cff_E[13] = 6'd2;                 assign ID_S_7f18c66f_6de04cff_E[14] = 6'd29;                 assign ID_S_7f18c66f_6de04cff_E[15] = 6'd28;             end          {4'd6,6'd32}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 6'd17;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 6'd21;                 assign ID_S_7f18c66f_6de04cff_E[2 ] = 6'd55;                 assign ID_S_7f18c66f_6de04cff_E[3 ] = 6'd14;                 assign ID_S_7f18c66f_6de04cff_E[4 ] = 6'd36;                 assign ID_S_7f18c66f_6de04cff_E[5 ] = 6'd13;                 assign ID_S_7f18c66f_6de04cff_E[6 ] = 6'd27;                 assign ID_S_7f18c66f_6de04cff_E[7 ] = 6'd31;                 assign ID_S_7f18c66f_6de04cff_E[8 ] = 6'd62;                 assign ID_S_7f18c66f_6de04cff_E[9 ] = 6'd46;                 assign ID_S_7f18c66f_6de04cff_E[10] = 6'd26;                 assign ID_S_7f18c66f_6de04cff_E[11] = 6'd21;                 assign ID_S_7f18c66f_6de04cff_E[12] = 6'd12;                 assign ID_S_7f18c66f_6de04cff_E[13] = 6'd5;                 assign ID_S_7f18c66f_6de04cff_E[14] = 6'd57;                 assign ID_S_7f18c66f_6de04cff_E[15] = 6'd50;                 assign ID_S_7f18c66f_6de04cff_E[16] = 6'd55;                 assign ID_S_7f18c66f_6de04cff_E[17] = 6'd10;                 assign ID_S_7f18c66f_6de04cff_E[18] = 6'd62;                 assign ID_S_7f18c66f_6de04cff_E[19] = 6'd54;                 assign ID_S_7f18c66f_6de04cff_E[20] = 6'd4;                 assign ID_S_7f18c66f_6de04cff_E[21] = 6'd10;                 assign ID_S_7f18c66f_6de04cff_E[22] = 6'd47;                 assign ID_S_7f18c66f_6de04cff_E[23] = 6'd10;                 assign ID_S_7f18c66f_6de04cff_E[24] = 6'd25;                 assign ID_S_7f18c66f_6de04cff_E[25] = 6'd35;                 assign ID_S_7f18c66f_6de04cff_E[26] = 6'd41;                 assign ID_S_7f18c66f_6de04cff_E[27] = 6'd1;                 assign ID_S_7f18c66f_6de04cff_E[28] = 6'd19;                 assign ID_S_7f18c66f_6de04cff_E[29] = 6'd54;                 assign ID_S_7f18c66f_6de04cff_E[30] = 6'd53;                 assign ID_S_7f18c66f_6de04cff_E[31] = 6'd49;             end          {4'd7,6'd2}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 7'd8;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 7'd6;             end          {4'd7,6'd4}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 7'd72;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 7'd127;                 assign ID_S_7f18c66f_6de04cff_E[2 ] = 7'd81;                 assign ID_S_7f18c66f_6de04cff_E[3 ] = 7'd30;             end          {4'd7,6'd8}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 7'd96;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 7'd49;                 assign ID_S_7f18c66f_6de04cff_E[2 ] = 7'd62;                 assign ID_S_7f18c66f_6de04cff_E[3 ] = 7'd124;                 assign ID_S_7f18c66f_6de04cff_E[4 ] = 7'd64;                 assign ID_S_7f18c66f_6de04cff_E[5 ] = 7'd37;                 assign ID_S_7f18c66f_6de04cff_E[6 ] = 7'd24;                 assign ID_S_7f18c66f_6de04cff_E[7 ] = 7'd101;             end          {4'd7,6'd16}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 7'd36;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 7'd39;                 assign ID_S_7f18c66f_6de04cff_E[2 ] = 7'd10;                 assign ID_S_7f18c66f_6de04cff_E[3 ] = 7'd116;                 assign ID_S_7f18c66f_6de04cff_E[4 ] = 7'd4;                 assign ID_S_7f18c66f_6de04cff_E[5 ] = 7'd10;                 assign ID_S_7f18c66f_6de04cff_E[6 ] = 7'd122;                 assign ID_S_7f18c66f_6de04cff_E[7 ] = 7'd120;                 assign ID_S_7f18c66f_6de04cff_E[8 ] = 7'd72;                 assign ID_S_7f18c66f_6de04cff_E[9 ] = 7'd21;                 assign ID_S_7f18c66f_6de04cff_E[10] = 7'd27;                 assign ID_S_7f18c66f_6de04cff_E[11] = 7'd50;                 assign ID_S_7f18c66f_6de04cff_E[12] = 7'd70;                 assign ID_S_7f18c66f_6de04cff_E[13] = 7'd118;                 assign ID_S_7f18c66f_6de04cff_E[14] = 7'd89;                 assign ID_S_7f18c66f_6de04cff_E[15] = 7'd26;             end          {4'd7,6'd32}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 7'd114;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 7'd35;                 assign ID_S_7f18c66f_6de04cff_E[2 ] = 7'd60;                 assign ID_S_7f18c66f_6de04cff_E[3 ] = 7'd55;                 assign ID_S_7f18c66f_6de04cff_E[4 ] = 7'd32;                 assign ID_S_7f18c66f_6de04cff_E[5 ] = 7'd24;                 assign ID_S_7f18c66f_6de04cff_E[6 ] = 7'd63;                 assign ID_S_7f18c66f_6de04cff_E[7 ] = 7'd36;                 assign ID_S_7f18c66f_6de04cff_E[8 ] = 7'd87;                 assign ID_S_7f18c66f_6de04cff_E[9 ] = 7'd20;                 assign ID_S_7f18c66f_6de04cff_E[10] = 7'd77;                 assign ID_S_7f18c66f_6de04cff_E[11] = 7'd32;                 assign ID_S_7f18c66f_6de04cff_E[12] = 7'd76;                 assign ID_S_7f18c66f_6de04cff_E[13] = 7'd52;                 assign ID_S_7f18c66f_6de04cff_E[14] = 7'd108;                 assign ID_S_7f18c66f_6de04cff_E[15] = 7'd58;                 assign ID_S_7f18c66f_6de04cff_E[16] = 7'd126;                 assign ID_S_7f18c66f_6de04cff_E[17] = 7'd65;                 assign ID_S_7f18c66f_6de04cff_E[18] = 7'd103;                 assign ID_S_7f18c66f_6de04cff_E[19] = 7'd79;                 assign ID_S_7f18c66f_6de04cff_E[20] = 7'd49;                 assign ID_S_7f18c66f_6de04cff_E[21] = 7'd30;                 assign ID_S_7f18c66f_6de04cff_E[22] = 7'd97;                 assign ID_S_7f18c66f_6de04cff_E[23] = 7'd104;                 assign ID_S_7f18c66f_6de04cff_E[24] = 7'd80;                 assign ID_S_7f18c66f_6de04cff_E[25] = 7'd15;                 assign ID_S_7f18c66f_6de04cff_E[26] = 7'd24;                 assign ID_S_7f18c66f_6de04cff_E[27] = 7'd62;                 assign ID_S_7f18c66f_6de04cff_E[28] = 7'd92;                 assign ID_S_7f18c66f_6de04cff_E[29] = 7'd36;                 assign ID_S_7f18c66f_6de04cff_E[30] = 7'd65;                 assign ID_S_7f18c66f_6de04cff_E[31] = 7'd125;             end                              {4'd8,6'd2}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 8'd8;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 8'd6;             end          {4'd8,6'd4}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 8'd116;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 8'd231;                 assign ID_S_7f18c66f_6de04cff_E[2 ] = 8'd216;                 assign ID_S_7f18c66f_6de04cff_E[3 ] = 8'd30;             end          {4'd8,6'd8}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 8'd37;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 8'd224;                 assign ID_S_7f18c66f_6de04cff_E[2 ] = 8'd8;                 assign ID_S_7f18c66f_6de04cff_E[3 ] = 8'd172;                 assign ID_S_7f18c66f_6de04cff_E[4 ] = 8'd71;                 assign ID_S_7f18c66f_6de04cff_E[5 ] = 8'd178;                 assign ID_S_7f18c66f_6de04cff_E[6 ] = 8'd44;                 assign ID_S_7f18c66f_6de04cff_E[7 ] = 8'd227;             end          {4'd8,6'd16}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 8'd79;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 8'd44;                 assign ID_S_7f18c66f_6de04cff_E[2 ] = 8'd81;                 assign ID_S_7f18c66f_6de04cff_E[3 ] = 8'd100;                 assign ID_S_7f18c66f_6de04cff_E[4 ] = 8'd49;                 assign ID_S_7f18c66f_6de04cff_E[5 ] = 8'd183;                 assign ID_S_7f18c66f_6de04cff_E[6 ] = 8'd56;                 assign ID_S_7f18c66f_6de04cff_E[7 ] = 8'd17;                 assign ID_S_7f18c66f_6de04cff_E[8 ] = 8'd232;                 assign ID_S_7f18c66f_6de04cff_E[9 ] = 8'd187;                 assign ID_S_7f18c66f_6de04cff_E[10] = 8'd126;                 assign ID_S_7f18c66f_6de04cff_E[11] = 8'd104;                 assign ID_S_7f18c66f_6de04cff_E[12] = 8'd31;                 assign ID_S_7f18c66f_6de04cff_E[13] = 8'd103;                 assign ID_S_7f18c66f_6de04cff_E[14] = 8'd52;                 assign ID_S_7f18c66f_6de04cff_E[15] = 8'd118;             end          {4'd8,6'd32}:             begin                 assign ID_S_7f18c66f_6de04cff_E[0 ] = 8'd45;                 assign ID_S_7f18c66f_6de04cff_E[1 ] = 8'd216;                 assign ID_S_7f18c66f_6de04cff_E[2 ] = 8'd239;                 assign ID_S_7f18c66f_6de04cff_E[3 ] = 8'd24;                 assign ID_S_7f18c66f_6de04cff_E[4 ] = 8'd253;                 assign ID_S_7f18c66f_6de04cff_E[5 ] = 8'd104;                 assign ID_S_7f18c66f_6de04cff_E[6 ] = 8'd27;                 assign ID_S_7f18c66f_6de04cff_E[7 ] = 8'd40;                 assign ID_S_7f18c66f_6de04cff_E[8 ] = 8'd107;                 assign ID_S_7f18c66f_6de04cff_E[9 ] = 8'd50;                 assign ID_S_7f18c66f_6de04cff_E[10] = 8'd163;                 assign ID_S_7f18c66f_6de04cff_E[11] = 8'd210;                 assign ID_S_7f18c66f_6de04cff_E[12] = 8'd227;                 assign ID_S_7f18c66f_6de04cff_E[13] = 8'd134;                 assign ID_S_7f18c66f_6de04cff_E[14] = 8'd224;                 assign ID_S_7f18c66f_6de04cff_E[15] = 8'd158;                 assign ID_S_7f18c66f_6de04cff_E[16] = 8'd119;                 assign ID_S_7f18c66f_6de04cff_E[17] = 8'd13;                 assign ID_S_7f18c66f_6de04cff_E[18] = 8'd158;                 assign ID_S_7f18c66f_6de04cff_E[19] = 8'd1;                 assign ID_S_7f18c66f_6de04cff_E[20] = 8'd238;                 assign ID_S_7f18c66f_6de04cff_E[21] = 8'd164;                 assign ID_S_7f18c66f_6de04cff_E[22] = 8'd82;                 assign ID_S_7f18c66f_6de04cff_E[23] = 8'd43;                 assign ID_S_7f18c66f_6de04cff_E[24] = 8'd15;                 assign ID_S_7f18c66f_6de04cff_E[25] = 8'd232;                 assign ID_S_7f18c66f_6de04cff_E[26] = 8'd246;                 assign ID_S_7f18c66f_6de04cff_E[27] = 8'd142;                 assign ID_S_7f18c66f_6de04cff_E[28] = 8'd50;                 assign ID_S_7f18c66f_6de04cff_E[29] = 8'd189;                 assign ID_S_7f18c66f_6de04cff_E[30] = 8'd29;                 assign ID_S_7f18c66f_6de04cff_E[31] = 8'd232;             end                                     endcase endgenerate   reg  [SYM_BW-1 :0] ID_S_3f3f4165_4359b2fd_E;   always @(posedge clk or negedge rst_n) if (!rst_n)   ID_S_3f3f4165_4359b2fd_E <= 0;   else if(din_sop == 1)   ID_S_3f3f4165_4359b2fd_E <= 1; else if(ID_S_3f3f4165_4359b2fd_E != 0 && ID_S_3f3f4165_4359b2fd_E < N_NUM)   ID_S_3f3f4165_4359b2fd_E <= ID_S_3f3f4165_4359b2fd_E + 1;   else    ID_S_3f3f4165_4359b2fd_E <= 0;    reg   [SYM_BW-1:0] ID_S_601727a0_6102309f_E     [R_NUM - 1:0]; wire  [SYM_BW-1:0] ID_S_60d7f109_28c363d0_E [R_NUM - 1:0]; wire  [SYM_BW-1:0] ID_S_4337be46_63201458_E      [R_NUM - 1:0];   wire  [SYM_BW-1:0] ID_S_35292296_41a22a95_E     [R_NUM - 1:0]; wire  [SYM_BW-1:0] ID_S_13ba76ff_5a73b221_E [R_NUM - 1:0];    genvar ID_S_1043cd9b_63834a56_E; generate     for(ID_S_1043cd9b_63834a56_E = 0;ID_S_1043cd9b_63834a56_E < R_NUM ;ID_S_1043cd9b_63834a56_E = ID_S_1043cd9b_63834a56_E + 1)     begin         always @(posedge clk or negedge rst_n)         if (!rst_n) begin           ID_S_601727a0_6102309f_E[ID_S_1043cd9b_63834a56_E] <= 0;           end else begin           ID_S_601727a0_6102309f_E[ID_S_1043cd9b_63834a56_E] <= ID_S_60d7f109_28c363d0_E[ID_S_1043cd9b_63834a56_E];           end     end endgenerate    reg [SYM_BW-1:0] ID_S_60d7f757_28c7eb46_E; always @(posedge clk or negedge rst_n) if (!rst_n) begin   ID_S_60d7f757_28c7eb46_E <= 0;  end else begin   ID_S_60d7f757_28c7eb46_E <= ID_S_601727a0_6102309f_E[R_NUM - 1];  end       reg [SYM_BW-1:0] ID_S_f4c06e3_2b609816_E;   always @(posedge clk or negedge rst_n) if (!rst_n)   ID_S_f4c06e3_2b609816_E <= 0;   else   ID_S_f4c06e3_2b609816_E <= din;    wire [SYM_BW-1:0] ID_S_6096e3a9_407934b0_E;  assign   ID_S_6096e3a9_407934b0_E = (din_val)? (din ^ ID_S_601727a0_6102309f_E[R_NUM - 1] ): 0;        generate     for(ID_S_1043cd9b_63834a56_E = 0;ID_S_1043cd9b_63834a56_E < R_NUM ;ID_S_1043cd9b_63834a56_E = ID_S_1043cd9b_63834a56_E + 1)     begin         case({ID_S_12846e01_7d0ea1dd_E})             {4'd3}:             begin                 gf8mul ID_S_44f4845b_5a564e7c_E (ID_S_6096e3a9_407934b0_E, ID_S_7f18c66f_6de04cff_E[ID_S_1043cd9b_63834a56_E], ID_S_4337be46_63201458_E[ID_S_1043cd9b_63834a56_E]);                         end                         {4'd4}:             begin                 gf16mul ID_S_44f4845b_5a564e7c_E (ID_S_6096e3a9_407934b0_E, ID_S_7f18c66f_6de04cff_E[ID_S_1043cd9b_63834a56_E], ID_S_4337be46_63201458_E[ID_S_1043cd9b_63834a56_E]);                       end               {4'd5}:             begin                 gf32mul ID_S_44f4845b_5a564e7c_E (ID_S_6096e3a9_407934b0_E, ID_S_7f18c66f_6de04cff_E[ID_S_1043cd9b_63834a56_E], ID_S_4337be46_63201458_E[ID_S_1043cd9b_63834a56_E]);                       end                         {4'd6}:             begin                 gf64mul ID_S_44f4845b_5a564e7c_E (ID_S_6096e3a9_407934b0_E, ID_S_7f18c66f_6de04cff_E[ID_S_1043cd9b_63834a56_E], ID_S_4337be46_63201458_E[ID_S_1043cd9b_63834a56_E]);                        end                         {4'd7}:             begin                 gf128mul ID_S_44f4845b_5a564e7c_E (ID_S_6096e3a9_407934b0_E, ID_S_7f18c66f_6de04cff_E[ID_S_1043cd9b_63834a56_E], ID_S_4337be46_63201458_E[ID_S_1043cd9b_63834a56_E]);                         end                       {4'd8}:             begin                 gf256mul ID_S_44f4845b_5a564e7c_E (ID_S_6096e3a9_407934b0_E, ID_S_7f18c66f_6de04cff_E[ID_S_1043cd9b_63834a56_E], ID_S_4337be46_63201458_E[ID_S_1043cd9b_63834a56_E]);                         end         endcase                    end endgenerate    assign  ID_S_60d7f109_28c363d0_E[0] = ID_S_4337be46_63201458_E[0];   generate     for(ID_S_1043cd9b_63834a56_E = 1;ID_S_1043cd9b_63834a56_E < R_NUM ;ID_S_1043cd9b_63834a56_E = ID_S_1043cd9b_63834a56_E + 1)     begin         assign  ID_S_60d7f109_28c363d0_E[ID_S_1043cd9b_63834a56_E] = ID_S_4337be46_63201458_E[ID_S_1043cd9b_63834a56_E] ^ ID_S_601727a0_6102309f_E[ID_S_1043cd9b_63834a56_E - 1];     end endgenerate  always @(posedge clk or negedge rst_n) if (!rst_n) begin   dout <= 0;  end else if(ID_S_3f3f4165_4359b2fd_E <= (N_NUM - R_NUM) && ID_S_3f3f4165_4359b2fd_E != 0) begin   dout <= ID_S_f4c06e3_2b609816_E;  end else if(ID_S_3f3f4165_4359b2fd_E > (N_NUM - R_NUM) && ID_S_3f3f4165_4359b2fd_E <= N_NUM) begin   dout <= ID_S_60d7f757_28c7eb46_E;    end else   dout <= 0;       always @(posedge clk or negedge rst_n) if (!rst_n) begin   dout_val <= 0;  end else   dout_val <= (ID_S_3f3f4165_4359b2fd_E != 0) && (ID_S_3f3f4165_4359b2fd_E <= N_NUM);     always @(posedge clk or negedge rst_n) if (!rst_n) begin   dout_sop <= 0;  end else   dout_sop <= (ID_S_3f3f4165_4359b2fd_E == 1);     always @(posedge clk or negedge rst_n) if (!rst_n) begin   dout_eop <= 0;  end else   dout_eop <= (ID_S_3f3f4165_4359b2fd_E == N_NUM);   endmodule