`timescale 1ns/100ps
////////////////////////////////////////////////////////////////
module idx2gf8(
       input [2:0] idx,
       output reg [2:0] z
       );
                                                                             
always @( * ) begin
  case (idx) 
	3'd  0: z = 3'd1;   
	3'd  1: z = 3'd2;  //a^0
	3'd  2: z = 3'd4;  //a^1
	3'd  3: z = 3'd3;
	3'd  4: z = 3'd6;
	3'd  5: z = 3'd7;
	3'd  6: z = 3'd5;
	3'd  7: z = 3'd1;
endcase
end
endmodule

////////////////////////////////////////////////////////////////
module idx2gf16(
       input [3:0] idx,
       output reg [3:0] z
       );
                                                                             
always @( * ) begin
  case (idx) 
	4'd  0: z = 4'd 1;   
	4'd  1: z = 4'd 2;  //a^0
	4'd  2: z = 4'd 4;  //a^1
	4'd  3: z = 4'd 8;
	4'd  4: z = 4'd 3;
	4'd  5: z = 4'd 6;
	4'd  6: z = 4'd12;
	4'd  7: z = 4'd11;
	4'd  8: z = 4'd 5;
	4'd  9: z = 4'd10;
	4'd 10: z = 4'd 7;
	4'd 11: z = 4'd14;
	4'd 12: z = 4'd15;
	4'd 13: z = 4'd13;
	4'd 14: z = 4'd 9;
	4'd 15: z = 4'd 1;
endcase
end
endmodule


////////////////////////////////////////////////////////////////
module idx2gf32(
       input [4:0] idx,
       output reg [4:0] z
       );
                                                                             
always @( * ) begin
  case (idx) 
	5'd  0: z = 5'd 1;   
	5'd  1: z = 5'd 2;  //a^0
	5'd  2: z = 5'd 4;  //a^1
	5'd  3: z = 5'd 8;
	5'd  4: z = 5'd16;
	5'd  5: z = 5'd 5;
	5'd  6: z = 5'd10;
	5'd  7: z = 5'd20;
	5'd  8: z = 5'd13;
	5'd  9: z = 5'd26;
	5'd 10: z = 5'd17;
	5'd 11: z = 5'd 7;
	5'd 12: z = 5'd14;
	5'd 13: z = 5'd28;
	5'd 14: z = 5'd29;
	5'd 15: z = 5'd31;
	5'd 16: z = 5'd27;
	5'd 17: z = 5'd19;
	5'd 18: z = 5'd 3;
	5'd 19: z = 5'd 6;
	5'd 20: z = 5'd12;
	5'd 21: z = 5'd24;
	5'd 22: z = 5'd21;
	5'd 23: z = 5'd15;
	5'd 24: z = 5'd30;
	5'd 25: z = 5'd25;
	5'd 26: z = 5'd23;
	5'd 27: z = 5'd11;
	5'd 28: z = 5'd22;
	5'd 29: z = 5'd 9;
	5'd 30: z = 5'd18;
	5'd 31: z = 5'd 1;
endcase
end
endmodule
 
////////////////////////////////////////////////////////////////
module idx2gf64(
       input [5:0] idx,
       output reg [5:0] z
       );
                                                                             
always @( * ) begin
  case (idx) 
	6'd  0: z = 6'd  1;   
	6'd  1: z = 6'd  2;  //a^0
	6'd  2: z = 6'd  4;  //a^1
	6'd  3: z = 6'd  8;
	6'd  4: z = 6'd 16;
	6'd  5: z = 6'd 32;
	6'd  6: z = 6'd  3;
	6'd  7: z = 6'd  6;
	6'd  8: z = 6'd 12;
	6'd  9: z = 6'd 24;
	6'd 10: z = 6'd 48;
	6'd 11: z = 6'd 35;
	6'd 12: z = 6'd  5;
	6'd 13: z = 6'd 10;
	6'd 14: z = 6'd 20;
	6'd 15: z = 6'd 40;
	6'd 16: z = 6'd 19;
	6'd 17: z = 6'd 38;
	6'd 18: z = 6'd 15;
	6'd 19: z = 6'd 30;
	6'd 20: z = 6'd 60;
	6'd 21: z = 6'd 59;
	6'd 22: z = 6'd 53;
	6'd 23: z = 6'd 41;
	6'd 24: z = 6'd 17;
	6'd 25: z = 6'd 34;
	6'd 26: z = 6'd  7;
	6'd 27: z = 6'd 14;
	6'd 28: z = 6'd 28;
	6'd 29: z = 6'd 56;
	6'd 30: z = 6'd 51;
	6'd 31: z = 6'd 37;
	6'd 32: z = 6'd  9;
	6'd 33: z = 6'd 18;
	6'd 34: z = 6'd 36;
	6'd 35: z = 6'd 11;
	6'd 36: z = 6'd 22;
	6'd 37: z = 6'd 44;
	6'd 38: z = 6'd 27;
	6'd 39: z = 6'd 54;
	6'd 40: z = 6'd 47;
	6'd 41: z = 6'd 29;
	6'd 42: z = 6'd 58;
	6'd 43: z = 6'd 55;
	6'd 44: z = 6'd 45;
	6'd 45: z = 6'd 25;
	6'd 46: z = 6'd 50;
	6'd 47: z = 6'd 39;
	6'd 48: z = 6'd 13;
	6'd 49: z = 6'd 26;
	6'd 50: z = 6'd 52;
	6'd 51: z = 6'd 43;
	6'd 52: z = 6'd 21;
	6'd 53: z = 6'd 42;
	6'd 54: z = 6'd 23;
	6'd 55: z = 6'd 46;
	6'd 56: z = 6'd 31;
	6'd 57: z = 6'd 62;
	6'd 58: z = 6'd 63;
	6'd 59: z = 6'd 61;
	6'd 60: z = 6'd 57;
	6'd 61: z = 6'd 49;
	6'd 62: z = 6'd 33;
	6'd 63: z = 6'd  1;

endcase
end
endmodule

////////////////////////////////////////////////////////////////
module idx2gf128(
       input [6:0] idx,
       output reg [6:0] z
       );
                                                                             
always @( * ) begin
  case (idx) 
	7'd  0: z = 7'd  1;   
	7'd  1: z = 7'd  2;  //a^0
	7'd  2: z = 7'd  4;  //a^1
	7'd  3: z = 7'd  8;
	7'd  4: z = 7'd 16;
	7'd  5: z = 7'd 32;
	7'd  6: z = 7'd 64;
	7'd  7: z = 7'd  9;
	7'd  8: z = 7'd 18;
	7'd  9: z = 7'd 36;
	7'd 10: z = 7'd 72;
	7'd 11: z = 7'd 25;
	7'd 12: z = 7'd 50;
	7'd 13: z = 7'd100;
	7'd 14: z = 7'd 65;
	7'd 15: z = 7'd 11;
	7'd 16: z = 7'd 22;
	7'd 17: z = 7'd 44;
	7'd 18: z = 7'd 88;
	7'd 19: z = 7'd 57;
	7'd 20: z = 7'd114;
	7'd 21: z = 7'd109;
	7'd 22: z = 7'd 83;
	7'd 23: z = 7'd 47;
	7'd 24: z = 7'd 94;
	7'd 25: z = 7'd 53;
	7'd 26: z = 7'd106;
	7'd 27: z = 7'd 93;
	7'd 28: z = 7'd 51;
	7'd 29: z = 7'd102;
	7'd 30: z = 7'd 69;
	7'd 31: z = 7'd  3;
	7'd 32: z = 7'd  6;
	7'd 33: z = 7'd 12;
	7'd 34: z = 7'd 24;
	7'd 35: z = 7'd 48;
	7'd 36: z = 7'd 96;
	7'd 37: z = 7'd 73;
	7'd 38: z = 7'd 27;
	7'd 39: z = 7'd 54;
	7'd 40: z = 7'd108;
	7'd 41: z = 7'd 81;
	7'd 42: z = 7'd 43;
	7'd 43: z = 7'd 86;
	7'd 44: z = 7'd 37;
	7'd 45: z = 7'd 74;
	7'd 46: z = 7'd 29;
	7'd 47: z = 7'd 58;
	7'd 48: z = 7'd116;
	7'd 49: z = 7'd 97;
	7'd 50: z = 7'd 75;
	7'd 51: z = 7'd 31;
	7'd 52: z = 7'd 62;
	7'd 53: z = 7'd124;
	7'd 54: z = 7'd113;
	7'd 55: z = 7'd107;
	7'd 56: z = 7'd 95;
	7'd 57: z = 7'd 55;
	7'd 58: z = 7'd110;
	7'd 59: z = 7'd 85;
	7'd 60: z = 7'd 35;
	7'd 61: z = 7'd 70;
	7'd 62: z = 7'd  5;
	7'd 63: z = 7'd 10;
	7'd 64: z = 7'd 20;
	7'd 65: z = 7'd 40;
	7'd 66: z = 7'd 80;
	7'd 67: z = 7'd 41;
	7'd 68: z = 7'd 82;
	7'd 69: z = 7'd 45;
	7'd 70: z = 7'd 90;
	7'd 71: z = 7'd 61;
	7'd 72: z = 7'd122;
	7'd 73: z = 7'd125;
	7'd 74: z = 7'd115;
	7'd 75: z = 7'd111;
	7'd 76: z = 7'd 87;
	7'd 77: z = 7'd 39;
	7'd 78: z = 7'd 78;
	7'd 79: z = 7'd 21;
	7'd 80: z = 7'd 42;
	7'd 81: z = 7'd 84;
	7'd 82: z = 7'd 33;
	7'd 83: z = 7'd 66;
	7'd 84: z = 7'd 13;
	7'd 85: z = 7'd 26;
	7'd 86: z = 7'd 52;
	7'd 87: z = 7'd104;
	7'd 88: z = 7'd 89;
	7'd 89: z = 7'd 59;
	7'd 90: z = 7'd118;
	7'd 91: z = 7'd101;
	7'd 92: z = 7'd 67;
	7'd 93: z = 7'd 15;
	7'd 94: z = 7'd 30;
	7'd 95: z = 7'd 60;
	7'd 96: z = 7'd120;
	7'd 97: z = 7'd121;
	7'd 98: z = 7'd123;
	7'd 99: z = 7'd127;
	7'd100: z = 7'd119;
	7'd101: z = 7'd103;
	7'd102: z = 7'd 71;
	7'd103: z = 7'd  7;
	7'd104: z = 7'd 14;
	7'd105: z = 7'd 28;
	7'd106: z = 7'd 56;
	7'd107: z = 7'd112;
	7'd108: z = 7'd105;
	7'd109: z = 7'd 91;
	7'd110: z = 7'd 63;
	7'd111: z = 7'd126;
	7'd112: z = 7'd117;
	7'd113: z = 7'd 99;
	7'd114: z = 7'd 79;
	7'd115: z = 7'd 23;
	7'd116: z = 7'd 46;
	7'd117: z = 7'd 92;
	7'd118: z = 7'd 49;
	7'd119: z = 7'd 98;
	7'd120: z = 7'd 77;
	7'd121: z = 7'd 19;
	7'd122: z = 7'd 38;
	7'd123: z = 7'd 76;
	7'd124: z = 7'd 17;
	7'd125: z = 7'd 34;
	7'd126: z = 7'd 68;
	7'd127: z = 7'd  1;
endcase
end
endmodule
 


////////////////////////////////////////////////////////////////
module idx2gf256(
       input [7:0] idx,
       output reg [7:0] z
       );
                                                                             
always @( * ) begin
  case (idx) 
	8'd  0: z = 8'd  1;   
	8'd  1: z = 8'd  2;  //a^0
	8'd  2: z = 8'd  4;  //a^1
	8'd  3: z = 8'd  8;
	8'd  4: z = 8'd 16;
	8'd  5: z = 8'd 32;
	8'd  6: z = 8'd 64;
	8'd  7: z = 8'd128;
	8'd  8: z = 8'd 29;
	8'd  9: z = 8'd 58;
	8'd 10: z = 8'd116;
	8'd 11: z = 8'd232;
	8'd 12: z = 8'd205;
	8'd 13: z = 8'd135;
	8'd 14: z = 8'd 19;
	8'd 15: z = 8'd 38;
	8'd 16: z = 8'd 76;
	8'd 17: z = 8'd152;
	8'd 18: z = 8'd 45;
	8'd 19: z = 8'd 90;
	8'd 20: z = 8'd180;
	8'd 21: z = 8'd117;
	8'd 22: z = 8'd234;
	8'd 23: z = 8'd201;
	8'd 24: z = 8'd143;
	8'd 25: z = 8'd  3;
	8'd 26: z = 8'd  6;
	8'd 27: z = 8'd 12;
	8'd 28: z = 8'd 24;
	8'd 29: z = 8'd 48;
	8'd 30: z = 8'd 96;
	8'd 31: z = 8'd192;
	8'd 32: z = 8'd157;
	8'd 33: z = 8'd 39;
	8'd 34: z = 8'd 78;
	8'd 35: z = 8'd156;
	8'd 36: z = 8'd 37;
	8'd 37: z = 8'd 74;
	8'd 38: z = 8'd148;
	8'd 39: z = 8'd 53;
	8'd 40: z = 8'd106;
	8'd 41: z = 8'd212;
	8'd 42: z = 8'd181;
	8'd 43: z = 8'd119;
	8'd 44: z = 8'd238;
	8'd 45: z = 8'd193;
	8'd 46: z = 8'd159;
	8'd 47: z = 8'd 35;
	8'd 48: z = 8'd 70;
	8'd 49: z = 8'd140;
	8'd 50: z = 8'd  5;
	8'd 51: z = 8'd 10;
	8'd 52: z = 8'd 20;
	8'd 53: z = 8'd 40;
	8'd 54: z = 8'd 80;
	8'd 55: z = 8'd160;
	8'd 56: z = 8'd 93;
	8'd 57: z = 8'd186;
	8'd 58: z = 8'd105;
	8'd 59: z = 8'd210;
	8'd 60: z = 8'd185;
	8'd 61: z = 8'd111;
	8'd 62: z = 8'd222;
	8'd 63: z = 8'd161;
	8'd 64: z = 8'd 95;
	8'd 65: z = 8'd190;
	8'd 66: z = 8'd 97;
	8'd 67: z = 8'd194;
	8'd 68: z = 8'd153;
	8'd 69: z = 8'd 47;
	8'd 70: z = 8'd 94;
	8'd 71: z = 8'd188;
	8'd 72: z = 8'd101;
	8'd 73: z = 8'd202;
	8'd 74: z = 8'd137;
	8'd 75: z = 8'd 15;
	8'd 76: z = 8'd 30;
	8'd 77: z = 8'd 60;
	8'd 78: z = 8'd120;
	8'd 79: z = 8'd240;
	8'd 80: z = 8'd253;
	8'd 81: z = 8'd231;
	8'd 82: z = 8'd211;
	8'd 83: z = 8'd187;
	8'd 84: z = 8'd107;
	8'd 85: z = 8'd214;
	8'd 86: z = 8'd177;
	8'd 87: z = 8'd127;
	8'd 88: z = 8'd254;
	8'd 89: z = 8'd225;
	8'd 90: z = 8'd223;
	8'd 91: z = 8'd163;
	8'd 92: z = 8'd 91;
	8'd 93: z = 8'd182;
	8'd 94: z = 8'd113;
	8'd 95: z = 8'd226;
	8'd 96: z = 8'd217;
	8'd 97: z = 8'd175;
	8'd 98: z = 8'd 67;
	8'd 99: z = 8'd134;
	8'd100: z = 8'd 17;
	8'd101: z = 8'd 34;
	8'd102: z = 8'd 68;
	8'd103: z = 8'd136;
	8'd104: z = 8'd 13;
	8'd105: z = 8'd 26;
	8'd106: z = 8'd 52;
	8'd107: z = 8'd104;
	8'd108: z = 8'd208;
	8'd109: z = 8'd189;
	8'd110: z = 8'd103;
	8'd111: z = 8'd206;
	8'd112: z = 8'd129;
	8'd113: z = 8'd 31;
	8'd114: z = 8'd 62;
	8'd115: z = 8'd124;
	8'd116: z = 8'd248;
	8'd117: z = 8'd237;
	8'd118: z = 8'd199;
	8'd119: z = 8'd147;
	8'd120: z = 8'd 59;
	8'd121: z = 8'd118;
	8'd122: z = 8'd236;
	8'd123: z = 8'd197;
	8'd124: z = 8'd151;
	8'd125: z = 8'd 51;
	8'd126: z = 8'd102;
	8'd127: z = 8'd204;
	8'd128: z = 8'd133;
	8'd129: z = 8'd 23;
	8'd130: z = 8'd 46;
	8'd131: z = 8'd 92;
	8'd132: z = 8'd184;
	8'd133: z = 8'd109;
	8'd134: z = 8'd218;
	8'd135: z = 8'd169;
	8'd136: z = 8'd 79;
	8'd137: z = 8'd158;
	8'd138: z = 8'd 33;
	8'd139: z = 8'd 66;
	8'd140: z = 8'd132;
	8'd141: z = 8'd 21;
	8'd142: z = 8'd 42;
	8'd143: z = 8'd 84;
	8'd144: z = 8'd168;
	8'd145: z = 8'd 77;
	8'd146: z = 8'd154;
	8'd147: z = 8'd 41;
	8'd148: z = 8'd 82;
	8'd149: z = 8'd164;
	8'd150: z = 8'd 85;
	8'd151: z = 8'd170;
	8'd152: z = 8'd 73;
	8'd153: z = 8'd146;
	8'd154: z = 8'd 57;
	8'd155: z = 8'd114;
	8'd156: z = 8'd228;
	8'd157: z = 8'd213;
	8'd158: z = 8'd183;
	8'd159: z = 8'd115;
	8'd160: z = 8'd230;
	8'd161: z = 8'd209;
	8'd162: z = 8'd191;
	8'd163: z = 8'd 99;
	8'd164: z = 8'd198;
	8'd165: z = 8'd145;
	8'd166: z = 8'd 63;
	8'd167: z = 8'd126;
	8'd168: z = 8'd252;
	8'd169: z = 8'd229;
	8'd170: z = 8'd215;
	8'd171: z = 8'd179;
	8'd172: z = 8'd123;
	8'd173: z = 8'd246;
	8'd174: z = 8'd241;
	8'd175: z = 8'd255;
	8'd176: z = 8'd227;
	8'd177: z = 8'd219;
	8'd178: z = 8'd171;
	8'd179: z = 8'd 75;
	8'd180: z = 8'd150;
	8'd181: z = 8'd 49;
	8'd182: z = 8'd 98;
	8'd183: z = 8'd196;
	8'd184: z = 8'd149;
	8'd185: z = 8'd 55;
	8'd186: z = 8'd110;
	8'd187: z = 8'd220;
	8'd188: z = 8'd165;
	8'd189: z = 8'd 87;
	8'd190: z = 8'd174;
	8'd191: z = 8'd 65;
	8'd192: z = 8'd130;
	8'd193: z = 8'd 25;
	8'd194: z = 8'd 50;
	8'd195: z = 8'd100;
	8'd196: z = 8'd200;
	8'd197: z = 8'd141;
	8'd198: z = 8'd  7;
	8'd199: z = 8'd 14;
	8'd200: z = 8'd 28;
	8'd201: z = 8'd 56;
	8'd202: z = 8'd112;
	8'd203: z = 8'd224;
	8'd204: z = 8'd221;
	8'd205: z = 8'd167;
	8'd206: z = 8'd 83;
	8'd207: z = 8'd166;
	8'd208: z = 8'd 81;
	8'd209: z = 8'd162;
	8'd210: z = 8'd 89;
	8'd211: z = 8'd178;
	8'd212: z = 8'd121;
	8'd213: z = 8'd242;
	8'd214: z = 8'd249;
	8'd215: z = 8'd239;
	8'd216: z = 8'd195;
	8'd217: z = 8'd155;
	8'd218: z = 8'd 43;
	8'd219: z = 8'd 86;
	8'd220: z = 8'd172;
	8'd221: z = 8'd 69;
	8'd222: z = 8'd138;
	8'd223: z = 8'd  9;
	8'd224: z = 8'd 18;
	8'd225: z = 8'd 36;
	8'd226: z = 8'd 72;
	8'd227: z = 8'd144;
	8'd228: z = 8'd 61;
	8'd229: z = 8'd122;
	8'd230: z = 8'd244;
	8'd231: z = 8'd245;
	8'd232: z = 8'd247;
	8'd233: z = 8'd243;
	8'd234: z = 8'd251;
	8'd235: z = 8'd235;
	8'd236: z = 8'd203;
	8'd237: z = 8'd139;
	8'd238: z = 8'd 11;
	8'd239: z = 8'd 22;
	8'd240: z = 8'd 44;
	8'd241: z = 8'd 88;
	8'd242: z = 8'd176;
	8'd243: z = 8'd125;
	8'd244: z = 8'd250;
	8'd245: z = 8'd233;
	8'd246: z = 8'd207;
	8'd247: z = 8'd131;
	8'd248: z = 8'd 27;
	8'd249: z = 8'd 54;
	8'd250: z = 8'd108;
	8'd251: z = 8'd216;
	8'd252: z = 8'd173;
	8'd253: z = 8'd 71;
	8'd254: z = 8'd142;
	8'd255: z = 8'd1  ;
endcase
end


endmodule


